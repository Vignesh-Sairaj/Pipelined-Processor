`include "mux2to1.v"

`ifndef _Lshift24_
`define _Lshift24_

module Lshift24(A, shl, OUT);

	input [23:0] A;
	input [4:0] shl;

	output [23:0] OUT;

	wire [23:0] m0, m1, m2, m3, m4;

	reg z = 1'b0;

	mux2to1 M00(z, A[0], ~shl[0], m0[0]), M01(A[0], A[1], ~shl[0], m0[1]), M02(A[1], A[2], ~shl[0], m0[2]), M03(A[2], A[3], ~shl[0], m0[3]), M04(A[3], A[4], ~shl[0], m0[4]), M05(A[4], A[5], ~shl[0], m0[5]), M06(A[5], A[6], ~shl[0], m0[6]), M07(A[6], A[7], ~shl[0], m0[7]), M08(A[7], A[8], ~shl[0], m0[8]), M09(A[8], A[9], ~shl[0], m0[9]), M010(A[9], A[10], ~shl[0], m0[10]), M011(A[10], A[11], ~shl[0], m0[11]), M012(A[11], A[12], ~shl[0], m0[12]), M013(A[12], A[13], ~shl[0], m0[13]), M014(A[13], A[14], ~shl[0], m0[14]), M015(A[14], A[15], ~shl[0], m0[15]), M016(A[15], A[16], ~shl[0], m0[16]), M017(A[16], A[17], ~shl[0], m0[17]), M018(A[17], A[18], ~shl[0], m0[18]), M019(A[18], A[19], ~shl[0], m0[19]), M020(A[19], A[20], ~shl[0], m0[20]), M021(A[20], A[21], ~shl[0], m0[21]), M022(A[21], A[22], ~shl[0], m0[22]), M023(A[22], A[23], ~shl[0], m0[23]);

	mux2to1 M10(z, m0[0], ~shl[1], m1[0]), M11(z, m0[1], ~shl[1], m1[1]), M12(m0[0], m0[2], ~shl[1], m1[2]), M13(m0[1], m0[3], ~shl[1], m1[3]), M14(m0[2], m0[4], ~shl[1], m1[4]), M15(m0[3], m0[5], ~shl[1], m1[5]), M16(m0[4], m0[6], ~shl[1], m1[6]), M17(m0[5], m0[7], ~shl[1], m1[7]), M18(m0[6], m0[8], ~shl[1], m1[8]), M19(m0[7], m0[9], ~shl[1], m1[9]), M110(m0[8], m0[10], ~shl[1], m1[10]), M111(m0[9], m0[11], ~shl[1], m1[11]), M112(m0[10], m0[12], ~shl[1], m1[12]), M113(m0[11], m0[13], ~shl[1], m1[13]), M114(m0[12], m0[14], ~shl[1], m1[14]), M115(m0[13], m0[15], ~shl[1], m1[15]), M116(m0[14], m0[16], ~shl[1], m1[16]), M117(m0[15], m0[17], ~shl[1], m1[17]), M118(m0[16], m0[18], ~shl[1], m1[18]), M119(m0[17], m0[19], ~shl[1], m1[19]), M120(m0[18], m0[20], ~shl[1], m1[20]), M121(m0[19], m0[21], ~shl[1], m1[21]), M122(m0[20], m0[22], ~shl[1], m1[22]), M123(m0[21], m0[23], ~shl[1], m1[23]);

	mux2to1 M20(z, m1[0], ~shl[2], m2[0]), M21(z, m1[1], ~shl[2], m2[1]), M22(z, m1[2], ~shl[2], m2[2]), M23(z, m1[3], ~shl[2], m2[3]), M24(m1[0], m1[4], ~shl[2], m2[4]), M25(m1[1], m1[5], ~shl[2], m2[5]), M26(m1[2], m1[6], ~shl[2], m2[6]), M27(m1[3], m1[7], ~shl[2], m2[7]), M28(m1[4], m1[8], ~shl[2], m2[8]), M29(m1[5], m1[9], ~shl[2], m2[9]), M210(m1[6], m1[10], ~shl[2], m2[10]), M211(m1[7], m1[11], ~shl[2], m2[11]), M212(m1[8], m1[12], ~shl[2], m2[12]), M213(m1[9], m1[13], ~shl[2], m2[13]), M214(m1[10], m1[14], ~shl[2], m2[14]), M215(m1[11], m1[15], ~shl[2], m2[15]), M216(m1[12], m1[16], ~shl[2], m2[16]), M217(m1[13], m1[17], ~shl[2], m2[17]), M218(m1[14], m1[18], ~shl[2], m2[18]), M219(m1[15], m1[19], ~shl[2], m2[19]), M220(m1[16], m1[20], ~shl[2], m2[20]), M221(m1[17], m1[21], ~shl[2], m2[21]), M222(m1[18], m1[22], ~shl[2], m2[22]), M223(m1[19], m1[23], ~shl[2], m2[23]);

	mux2to1 M30(z, m2[0], ~shl[3], m3[0]), M31(z, m2[1], ~shl[3], m3[1]), M32(z, m2[2], ~shl[3], m3[2]), M33(z, m2[3], ~shl[3], m3[3]), M34(z, m2[4], ~shl[3], m3[4]), M35(z, m2[5], ~shl[3], m3[5]), M36(z, m2[6], ~shl[3], m3[6]), M37(z, m2[7], ~shl[3], m3[7]), M38(m2[0], m2[8], ~shl[3], m3[8]), M39(m2[1], m2[9], ~shl[3], m3[9]), M310(m2[2], m2[10], ~shl[3], m3[10]), M311(m2[3], m2[11], ~shl[3], m3[11]), M312(m2[4], m2[12], ~shl[3], m3[12]), M313(m2[5], m2[13], ~shl[3], m3[13]), M314(m2[6], m2[14], ~shl[3], m3[14]), M315(m2[7], m2[15], ~shl[3], m3[15]), M316(m2[8], m2[16], ~shl[3], m3[16]), M317(m2[9], m2[17], ~shl[3], m3[17]), M318(m2[10], m2[18], ~shl[3], m3[18]), M319(m2[11], m2[19], ~shl[3], m3[19]), M320(m2[12], m2[20], ~shl[3], m3[20]), M321(m2[13], m2[21], ~shl[3], m3[21]), M322(m2[14], m2[22], ~shl[3], m3[22]), M323(m2[15], m2[23], ~shl[3], m3[23]);

	mux2to1 M40(z, m3[0], ~shl[4], m4[0]), M41(z, m3[1], ~shl[4], m4[1]), M42(z, m3[2], ~shl[4], m4[2]), M43(z, m3[3], ~shl[4], m4[3]), M44(z, m3[4], ~shl[4], m4[4]), M45(z, m3[5], ~shl[4], m4[5]), M46(z, m3[6], ~shl[4], m4[6]), M47(z, m3[7], ~shl[4], m4[7]), M48(z, m3[8], ~shl[4], m4[8]), M49(z, m3[9], ~shl[4], m4[9]), M410(z, m3[10], ~shl[4], m4[10]), M411(z, m3[11], ~shl[4], m4[11]), M412(z, m3[12], ~shl[4], m4[12]), M413(z, m3[13], ~shl[4], m4[13]), M414(z, m3[14], ~shl[4], m4[14]), M415(z, m3[15], ~shl[4], m4[15]), M416(m3[0], m3[16], ~shl[4], m4[16]), M417(m3[1], m3[17], ~shl[4], m4[17]), M418(m3[2], m3[18], ~shl[4], m4[18]), M419(m3[3], m3[19], ~shl[4], m4[19]), M420(m3[4], m3[20], ~shl[4], m4[20]), M421(m3[5], m3[21], ~shl[4], m4[21]), M422(m3[6], m3[22], ~shl[4], m4[22]), M423(m3[7], m3[23], ~shl[4], m4[23]);

	assign OUT = m4;
endmodule
`endif