module CLA_48(x, y, cIn, s, cOut);

	input [47:0] x, y;
	input cIn;

	output [47:0] s;
	output cOut;

	wire [47:0] g, p;
	wire [48:0] c;

	assign g = x&y;
	assign p = x^y;

	assign c[0] = cIn;

	assign c[1] = g[0] | &p[0:0]&c[0];
	assign c[2] = g[1] | &p[1:1]&g[0] | &p[1:0]&c[0];
	assign c[3] = g[2] | &p[2:2]&g[1] | &p[2:1]&g[0] | &p[2:0]&c[0];
	assign c[4] = g[3] | &p[3:3]&g[2] | &p[3:2]&g[1] | &p[3:1]&g[0] | &p[3:0]&c[0];
	assign c[5] = g[4] | &p[4:4]&g[3] | &p[4:3]&g[2] | &p[4:2]&g[1] | &p[4:1]&g[0] | &p[4:0]&c[0];
	assign c[6] = g[5] | &p[5:5]&g[4] | &p[5:4]&g[3] | &p[5:3]&g[2] | &p[5:2]&g[1] | &p[5:1]&g[0] | &p[5:0]&c[0];
	assign c[7] = g[6] | &p[6:6]&g[5] | &p[6:5]&g[4] | &p[6:4]&g[3] | &p[6:3]&g[2] | &p[6:2]&g[1] | &p[6:1]&g[0] | &p[6:0]&c[0];
	assign c[8] = g[7] | &p[7:7]&g[6] | &p[7:6]&g[5] | &p[7:5]&g[4] | &p[7:4]&g[3] | &p[7:3]&g[2] | &p[7:2]&g[1] | &p[7:1]&g[0] | &p[7:0]&c[0];
	assign c[9] = g[8] | &p[8:8]&g[7] | &p[8:7]&g[6] | &p[8:6]&g[5] | &p[8:5]&g[4] | &p[8:4]&g[3] | &p[8:3]&g[2] | &p[8:2]&g[1] | &p[8:1]&g[0] | &p[8:0]&c[0];
	assign c[10] = g[9] | &p[9:9]&g[8] | &p[9:8]&g[7] | &p[9:7]&g[6] | &p[9:6]&g[5] | &p[9:5]&g[4] | &p[9:4]&g[3] | &p[9:3]&g[2] | &p[9:2]&g[1] | &p[9:1]&g[0] | &p[9:0]&c[0];
	assign c[11] = g[10] | &p[10:10]&g[9] | &p[10:9]&g[8] | &p[10:8]&g[7] | &p[10:7]&g[6] | &p[10:6]&g[5] | &p[10:5]&g[4] | &p[10:4]&g[3] | &p[10:3]&g[2] | &p[10:2]&g[1] | &p[10:1]&g[0] | &p[10:0]&c[0];
	assign c[12] = g[11] | &p[11:11]&g[10] | &p[11:10]&g[9] | &p[11:9]&g[8] | &p[11:8]&g[7] | &p[11:7]&g[6] | &p[11:6]&g[5] | &p[11:5]&g[4] | &p[11:4]&g[3] | &p[11:3]&g[2] | &p[11:2]&g[1] | &p[11:1]&g[0] | &p[11:0]&c[0];
	assign c[13] = g[12] | &p[12:12]&g[11] | &p[12:11]&g[10] | &p[12:10]&g[9] | &p[12:9]&g[8] | &p[12:8]&g[7] | &p[12:7]&g[6] | &p[12:6]&g[5] | &p[12:5]&g[4] | &p[12:4]&g[3] | &p[12:3]&g[2] | &p[12:2]&g[1] | &p[12:1]&g[0] | &p[12:0]&c[0];
	assign c[14] = g[13] | &p[13:13]&g[12] | &p[13:12]&g[11] | &p[13:11]&g[10] | &p[13:10]&g[9] | &p[13:9]&g[8] | &p[13:8]&g[7] | &p[13:7]&g[6] | &p[13:6]&g[5] | &p[13:5]&g[4] | &p[13:4]&g[3] | &p[13:3]&g[2] | &p[13:2]&g[1] | &p[13:1]&g[0] | &p[13:0]&c[0];
	assign c[15] = g[14] | &p[14:14]&g[13] | &p[14:13]&g[12] | &p[14:12]&g[11] | &p[14:11]&g[10] | &p[14:10]&g[9] | &p[14:9]&g[8] | &p[14:8]&g[7] | &p[14:7]&g[6] | &p[14:6]&g[5] | &p[14:5]&g[4] | &p[14:4]&g[3] | &p[14:3]&g[2] | &p[14:2]&g[1] | &p[14:1]&g[0] | &p[14:0]&c[0];
	assign c[16] = g[15] | &p[15:15]&g[14] | &p[15:14]&g[13] | &p[15:13]&g[12] | &p[15:12]&g[11] | &p[15:11]&g[10] | &p[15:10]&g[9] | &p[15:9]&g[8] | &p[15:8]&g[7] | &p[15:7]&g[6] | &p[15:6]&g[5] | &p[15:5]&g[4] | &p[15:4]&g[3] | &p[15:3]&g[2] | &p[15:2]&g[1] | &p[15:1]&g[0] | &p[15:0]&c[0];
	assign c[17] = g[16] | &p[16:16]&g[15] | &p[16:15]&g[14] | &p[16:14]&g[13] | &p[16:13]&g[12] | &p[16:12]&g[11] | &p[16:11]&g[10] | &p[16:10]&g[9] | &p[16:9]&g[8] | &p[16:8]&g[7] | &p[16:7]&g[6] | &p[16:6]&g[5] | &p[16:5]&g[4] | &p[16:4]&g[3] | &p[16:3]&g[2] | &p[16:2]&g[1] | &p[16:1]&g[0] | &p[16:0]&c[0];
	assign c[18] = g[17] | &p[17:17]&g[16] | &p[17:16]&g[15] | &p[17:15]&g[14] | &p[17:14]&g[13] | &p[17:13]&g[12] | &p[17:12]&g[11] | &p[17:11]&g[10] | &p[17:10]&g[9] | &p[17:9]&g[8] | &p[17:8]&g[7] | &p[17:7]&g[6] | &p[17:6]&g[5] | &p[17:5]&g[4] | &p[17:4]&g[3] | &p[17:3]&g[2] | &p[17:2]&g[1] | &p[17:1]&g[0] | &p[17:0]&c[0];
	assign c[19] = g[18] | &p[18:18]&g[17] | &p[18:17]&g[16] | &p[18:16]&g[15] | &p[18:15]&g[14] | &p[18:14]&g[13] | &p[18:13]&g[12] | &p[18:12]&g[11] | &p[18:11]&g[10] | &p[18:10]&g[9] | &p[18:9]&g[8] | &p[18:8]&g[7] | &p[18:7]&g[6] | &p[18:6]&g[5] | &p[18:5]&g[4] | &p[18:4]&g[3] | &p[18:3]&g[2] | &p[18:2]&g[1] | &p[18:1]&g[0] | &p[18:0]&c[0];
	assign c[20] = g[19] | &p[19:19]&g[18] | &p[19:18]&g[17] | &p[19:17]&g[16] | &p[19:16]&g[15] | &p[19:15]&g[14] | &p[19:14]&g[13] | &p[19:13]&g[12] | &p[19:12]&g[11] | &p[19:11]&g[10] | &p[19:10]&g[9] | &p[19:9]&g[8] | &p[19:8]&g[7] | &p[19:7]&g[6] | &p[19:6]&g[5] | &p[19:5]&g[4] | &p[19:4]&g[3] | &p[19:3]&g[2] | &p[19:2]&g[1] | &p[19:1]&g[0] | &p[19:0]&c[0];
	assign c[21] = g[20] | &p[20:20]&g[19] | &p[20:19]&g[18] | &p[20:18]&g[17] | &p[20:17]&g[16] | &p[20:16]&g[15] | &p[20:15]&g[14] | &p[20:14]&g[13] | &p[20:13]&g[12] | &p[20:12]&g[11] | &p[20:11]&g[10] | &p[20:10]&g[9] | &p[20:9]&g[8] | &p[20:8]&g[7] | &p[20:7]&g[6] | &p[20:6]&g[5] | &p[20:5]&g[4] | &p[20:4]&g[3] | &p[20:3]&g[2] | &p[20:2]&g[1] | &p[20:1]&g[0] | &p[20:0]&c[0];
	assign c[22] = g[21] | &p[21:21]&g[20] | &p[21:20]&g[19] | &p[21:19]&g[18] | &p[21:18]&g[17] | &p[21:17]&g[16] | &p[21:16]&g[15] | &p[21:15]&g[14] | &p[21:14]&g[13] | &p[21:13]&g[12] | &p[21:12]&g[11] | &p[21:11]&g[10] | &p[21:10]&g[9] | &p[21:9]&g[8] | &p[21:8]&g[7] | &p[21:7]&g[6] | &p[21:6]&g[5] | &p[21:5]&g[4] | &p[21:4]&g[3] | &p[21:3]&g[2] | &p[21:2]&g[1] | &p[21:1]&g[0] | &p[21:0]&c[0];
	assign c[23] = g[22] | &p[22:22]&g[21] | &p[22:21]&g[20] | &p[22:20]&g[19] | &p[22:19]&g[18] | &p[22:18]&g[17] | &p[22:17]&g[16] | &p[22:16]&g[15] | &p[22:15]&g[14] | &p[22:14]&g[13] | &p[22:13]&g[12] | &p[22:12]&g[11] | &p[22:11]&g[10] | &p[22:10]&g[9] | &p[22:9]&g[8] | &p[22:8]&g[7] | &p[22:7]&g[6] | &p[22:6]&g[5] | &p[22:5]&g[4] | &p[22:4]&g[3] | &p[22:3]&g[2] | &p[22:2]&g[1] | &p[22:1]&g[0] | &p[22:0]&c[0];
	assign c[24] = g[23] | &p[23:23]&g[22] | &p[23:22]&g[21] | &p[23:21]&g[20] | &p[23:20]&g[19] | &p[23:19]&g[18] | &p[23:18]&g[17] | &p[23:17]&g[16] | &p[23:16]&g[15] | &p[23:15]&g[14] | &p[23:14]&g[13] | &p[23:13]&g[12] | &p[23:12]&g[11] | &p[23:11]&g[10] | &p[23:10]&g[9] | &p[23:9]&g[8] | &p[23:8]&g[7] | &p[23:7]&g[6] | &p[23:6]&g[5] | &p[23:5]&g[4] | &p[23:4]&g[3] | &p[23:3]&g[2] | &p[23:2]&g[1] | &p[23:1]&g[0] | &p[23:0]&c[0];
	assign c[25] = g[24] | &p[24:24]&g[23] | &p[24:23]&g[22] | &p[24:22]&g[21] | &p[24:21]&g[20] | &p[24:20]&g[19] | &p[24:19]&g[18] | &p[24:18]&g[17] | &p[24:17]&g[16] | &p[24:16]&g[15] | &p[24:15]&g[14] | &p[24:14]&g[13] | &p[24:13]&g[12] | &p[24:12]&g[11] | &p[24:11]&g[10] | &p[24:10]&g[9] | &p[24:9]&g[8] | &p[24:8]&g[7] | &p[24:7]&g[6] | &p[24:6]&g[5] | &p[24:5]&g[4] | &p[24:4]&g[3] | &p[24:3]&g[2] | &p[24:2]&g[1] | &p[24:1]&g[0] | &p[24:0]&c[0];
	assign c[26] = g[25] | &p[25:25]&g[24] | &p[25:24]&g[23] | &p[25:23]&g[22] | &p[25:22]&g[21] | &p[25:21]&g[20] | &p[25:20]&g[19] | &p[25:19]&g[18] | &p[25:18]&g[17] | &p[25:17]&g[16] | &p[25:16]&g[15] | &p[25:15]&g[14] | &p[25:14]&g[13] | &p[25:13]&g[12] | &p[25:12]&g[11] | &p[25:11]&g[10] | &p[25:10]&g[9] | &p[25:9]&g[8] | &p[25:8]&g[7] | &p[25:7]&g[6] | &p[25:6]&g[5] | &p[25:5]&g[4] | &p[25:4]&g[3] | &p[25:3]&g[2] | &p[25:2]&g[1] | &p[25:1]&g[0] | &p[25:0]&c[0];
	assign c[27] = g[26] | &p[26:26]&g[25] | &p[26:25]&g[24] | &p[26:24]&g[23] | &p[26:23]&g[22] | &p[26:22]&g[21] | &p[26:21]&g[20] | &p[26:20]&g[19] | &p[26:19]&g[18] | &p[26:18]&g[17] | &p[26:17]&g[16] | &p[26:16]&g[15] | &p[26:15]&g[14] | &p[26:14]&g[13] | &p[26:13]&g[12] | &p[26:12]&g[11] | &p[26:11]&g[10] | &p[26:10]&g[9] | &p[26:9]&g[8] | &p[26:8]&g[7] | &p[26:7]&g[6] | &p[26:6]&g[5] | &p[26:5]&g[4] | &p[26:4]&g[3] | &p[26:3]&g[2] | &p[26:2]&g[1] | &p[26:1]&g[0] | &p[26:0]&c[0];
	assign c[28] = g[27] | &p[27:27]&g[26] | &p[27:26]&g[25] | &p[27:25]&g[24] | &p[27:24]&g[23] | &p[27:23]&g[22] | &p[27:22]&g[21] | &p[27:21]&g[20] | &p[27:20]&g[19] | &p[27:19]&g[18] | &p[27:18]&g[17] | &p[27:17]&g[16] | &p[27:16]&g[15] | &p[27:15]&g[14] | &p[27:14]&g[13] | &p[27:13]&g[12] | &p[27:12]&g[11] | &p[27:11]&g[10] | &p[27:10]&g[9] | &p[27:9]&g[8] | &p[27:8]&g[7] | &p[27:7]&g[6] | &p[27:6]&g[5] | &p[27:5]&g[4] | &p[27:4]&g[3] | &p[27:3]&g[2] | &p[27:2]&g[1] | &p[27:1]&g[0] | &p[27:0]&c[0];
	assign c[29] = g[28] | &p[28:28]&g[27] | &p[28:27]&g[26] | &p[28:26]&g[25] | &p[28:25]&g[24] | &p[28:24]&g[23] | &p[28:23]&g[22] | &p[28:22]&g[21] | &p[28:21]&g[20] | &p[28:20]&g[19] | &p[28:19]&g[18] | &p[28:18]&g[17] | &p[28:17]&g[16] | &p[28:16]&g[15] | &p[28:15]&g[14] | &p[28:14]&g[13] | &p[28:13]&g[12] | &p[28:12]&g[11] | &p[28:11]&g[10] | &p[28:10]&g[9] | &p[28:9]&g[8] | &p[28:8]&g[7] | &p[28:7]&g[6] | &p[28:6]&g[5] | &p[28:5]&g[4] | &p[28:4]&g[3] | &p[28:3]&g[2] | &p[28:2]&g[1] | &p[28:1]&g[0] | &p[28:0]&c[0];
	assign c[30] = g[29] | &p[29:29]&g[28] | &p[29:28]&g[27] | &p[29:27]&g[26] | &p[29:26]&g[25] | &p[29:25]&g[24] | &p[29:24]&g[23] | &p[29:23]&g[22] | &p[29:22]&g[21] | &p[29:21]&g[20] | &p[29:20]&g[19] | &p[29:19]&g[18] | &p[29:18]&g[17] | &p[29:17]&g[16] | &p[29:16]&g[15] | &p[29:15]&g[14] | &p[29:14]&g[13] | &p[29:13]&g[12] | &p[29:12]&g[11] | &p[29:11]&g[10] | &p[29:10]&g[9] | &p[29:9]&g[8] | &p[29:8]&g[7] | &p[29:7]&g[6] | &p[29:6]&g[5] | &p[29:5]&g[4] | &p[29:4]&g[3] | &p[29:3]&g[2] | &p[29:2]&g[1] | &p[29:1]&g[0] | &p[29:0]&c[0];
	assign c[31] = g[30] | &p[30:30]&g[29] | &p[30:29]&g[28] | &p[30:28]&g[27] | &p[30:27]&g[26] | &p[30:26]&g[25] | &p[30:25]&g[24] | &p[30:24]&g[23] | &p[30:23]&g[22] | &p[30:22]&g[21] | &p[30:21]&g[20] | &p[30:20]&g[19] | &p[30:19]&g[18] | &p[30:18]&g[17] | &p[30:17]&g[16] | &p[30:16]&g[15] | &p[30:15]&g[14] | &p[30:14]&g[13] | &p[30:13]&g[12] | &p[30:12]&g[11] | &p[30:11]&g[10] | &p[30:10]&g[9] | &p[30:9]&g[8] | &p[30:8]&g[7] | &p[30:7]&g[6] | &p[30:6]&g[5] | &p[30:5]&g[4] | &p[30:4]&g[3] | &p[30:3]&g[2] | &p[30:2]&g[1] | &p[30:1]&g[0] | &p[30:0]&c[0];
	assign c[32] = g[31] | &p[31:31]&g[30] | &p[31:30]&g[29] | &p[31:29]&g[28] | &p[31:28]&g[27] | &p[31:27]&g[26] | &p[31:26]&g[25] | &p[31:25]&g[24] | &p[31:24]&g[23] | &p[31:23]&g[22] | &p[31:22]&g[21] | &p[31:21]&g[20] | &p[31:20]&g[19] | &p[31:19]&g[18] | &p[31:18]&g[17] | &p[31:17]&g[16] | &p[31:16]&g[15] | &p[31:15]&g[14] | &p[31:14]&g[13] | &p[31:13]&g[12] | &p[31:12]&g[11] | &p[31:11]&g[10] | &p[31:10]&g[9] | &p[31:9]&g[8] | &p[31:8]&g[7] | &p[31:7]&g[6] | &p[31:6]&g[5] | &p[31:5]&g[4] | &p[31:4]&g[3] | &p[31:3]&g[2] | &p[31:2]&g[1] | &p[31:1]&g[0] | &p[31:0]&c[0];
	assign c[33] = g[32] | &p[32:32]&g[31] | &p[32:31]&g[30] | &p[32:30]&g[29] | &p[32:29]&g[28] | &p[32:28]&g[27] | &p[32:27]&g[26] | &p[32:26]&g[25] | &p[32:25]&g[24] | &p[32:24]&g[23] | &p[32:23]&g[22] | &p[32:22]&g[21] | &p[32:21]&g[20] | &p[32:20]&g[19] | &p[32:19]&g[18] | &p[32:18]&g[17] | &p[32:17]&g[16] | &p[32:16]&g[15] | &p[32:15]&g[14] | &p[32:14]&g[13] | &p[32:13]&g[12] | &p[32:12]&g[11] | &p[32:11]&g[10] | &p[32:10]&g[9] | &p[32:9]&g[8] | &p[32:8]&g[7] | &p[32:7]&g[6] | &p[32:6]&g[5] | &p[32:5]&g[4] | &p[32:4]&g[3] | &p[32:3]&g[2] | &p[32:2]&g[1] | &p[32:1]&g[0] | &p[32:0]&c[0];
	assign c[34] = g[33] | &p[33:33]&g[32] | &p[33:32]&g[31] | &p[33:31]&g[30] | &p[33:30]&g[29] | &p[33:29]&g[28] | &p[33:28]&g[27] | &p[33:27]&g[26] | &p[33:26]&g[25] | &p[33:25]&g[24] | &p[33:24]&g[23] | &p[33:23]&g[22] | &p[33:22]&g[21] | &p[33:21]&g[20] | &p[33:20]&g[19] | &p[33:19]&g[18] | &p[33:18]&g[17] | &p[33:17]&g[16] | &p[33:16]&g[15] | &p[33:15]&g[14] | &p[33:14]&g[13] | &p[33:13]&g[12] | &p[33:12]&g[11] | &p[33:11]&g[10] | &p[33:10]&g[9] | &p[33:9]&g[8] | &p[33:8]&g[7] | &p[33:7]&g[6] | &p[33:6]&g[5] | &p[33:5]&g[4] | &p[33:4]&g[3] | &p[33:3]&g[2] | &p[33:2]&g[1] | &p[33:1]&g[0] | &p[33:0]&c[0];
	assign c[35] = g[34] | &p[34:34]&g[33] | &p[34:33]&g[32] | &p[34:32]&g[31] | &p[34:31]&g[30] | &p[34:30]&g[29] | &p[34:29]&g[28] | &p[34:28]&g[27] | &p[34:27]&g[26] | &p[34:26]&g[25] | &p[34:25]&g[24] | &p[34:24]&g[23] | &p[34:23]&g[22] | &p[34:22]&g[21] | &p[34:21]&g[20] | &p[34:20]&g[19] | &p[34:19]&g[18] | &p[34:18]&g[17] | &p[34:17]&g[16] | &p[34:16]&g[15] | &p[34:15]&g[14] | &p[34:14]&g[13] | &p[34:13]&g[12] | &p[34:12]&g[11] | &p[34:11]&g[10] | &p[34:10]&g[9] | &p[34:9]&g[8] | &p[34:8]&g[7] | &p[34:7]&g[6] | &p[34:6]&g[5] | &p[34:5]&g[4] | &p[34:4]&g[3] | &p[34:3]&g[2] | &p[34:2]&g[1] | &p[34:1]&g[0] | &p[34:0]&c[0];
	assign c[36] = g[35] | &p[35:35]&g[34] | &p[35:34]&g[33] | &p[35:33]&g[32] | &p[35:32]&g[31] | &p[35:31]&g[30] | &p[35:30]&g[29] | &p[35:29]&g[28] | &p[35:28]&g[27] | &p[35:27]&g[26] | &p[35:26]&g[25] | &p[35:25]&g[24] | &p[35:24]&g[23] | &p[35:23]&g[22] | &p[35:22]&g[21] | &p[35:21]&g[20] | &p[35:20]&g[19] | &p[35:19]&g[18] | &p[35:18]&g[17] | &p[35:17]&g[16] | &p[35:16]&g[15] | &p[35:15]&g[14] | &p[35:14]&g[13] | &p[35:13]&g[12] | &p[35:12]&g[11] | &p[35:11]&g[10] | &p[35:10]&g[9] | &p[35:9]&g[8] | &p[35:8]&g[7] | &p[35:7]&g[6] | &p[35:6]&g[5] | &p[35:5]&g[4] | &p[35:4]&g[3] | &p[35:3]&g[2] | &p[35:2]&g[1] | &p[35:1]&g[0] | &p[35:0]&c[0];
	assign c[37] = g[36] | &p[36:36]&g[35] | &p[36:35]&g[34] | &p[36:34]&g[33] | &p[36:33]&g[32] | &p[36:32]&g[31] | &p[36:31]&g[30] | &p[36:30]&g[29] | &p[36:29]&g[28] | &p[36:28]&g[27] | &p[36:27]&g[26] | &p[36:26]&g[25] | &p[36:25]&g[24] | &p[36:24]&g[23] | &p[36:23]&g[22] | &p[36:22]&g[21] | &p[36:21]&g[20] | &p[36:20]&g[19] | &p[36:19]&g[18] | &p[36:18]&g[17] | &p[36:17]&g[16] | &p[36:16]&g[15] | &p[36:15]&g[14] | &p[36:14]&g[13] | &p[36:13]&g[12] | &p[36:12]&g[11] | &p[36:11]&g[10] | &p[36:10]&g[9] | &p[36:9]&g[8] | &p[36:8]&g[7] | &p[36:7]&g[6] | &p[36:6]&g[5] | &p[36:5]&g[4] | &p[36:4]&g[3] | &p[36:3]&g[2] | &p[36:2]&g[1] | &p[36:1]&g[0] | &p[36:0]&c[0];
	assign c[38] = g[37] | &p[37:37]&g[36] | &p[37:36]&g[35] | &p[37:35]&g[34] | &p[37:34]&g[33] | &p[37:33]&g[32] | &p[37:32]&g[31] | &p[37:31]&g[30] | &p[37:30]&g[29] | &p[37:29]&g[28] | &p[37:28]&g[27] | &p[37:27]&g[26] | &p[37:26]&g[25] | &p[37:25]&g[24] | &p[37:24]&g[23] | &p[37:23]&g[22] | &p[37:22]&g[21] | &p[37:21]&g[20] | &p[37:20]&g[19] | &p[37:19]&g[18] | &p[37:18]&g[17] | &p[37:17]&g[16] | &p[37:16]&g[15] | &p[37:15]&g[14] | &p[37:14]&g[13] | &p[37:13]&g[12] | &p[37:12]&g[11] | &p[37:11]&g[10] | &p[37:10]&g[9] | &p[37:9]&g[8] | &p[37:8]&g[7] | &p[37:7]&g[6] | &p[37:6]&g[5] | &p[37:5]&g[4] | &p[37:4]&g[3] | &p[37:3]&g[2] | &p[37:2]&g[1] | &p[37:1]&g[0] | &p[37:0]&c[0];
	assign c[39] = g[38] | &p[38:38]&g[37] | &p[38:37]&g[36] | &p[38:36]&g[35] | &p[38:35]&g[34] | &p[38:34]&g[33] | &p[38:33]&g[32] | &p[38:32]&g[31] | &p[38:31]&g[30] | &p[38:30]&g[29] | &p[38:29]&g[28] | &p[38:28]&g[27] | &p[38:27]&g[26] | &p[38:26]&g[25] | &p[38:25]&g[24] | &p[38:24]&g[23] | &p[38:23]&g[22] | &p[38:22]&g[21] | &p[38:21]&g[20] | &p[38:20]&g[19] | &p[38:19]&g[18] | &p[38:18]&g[17] | &p[38:17]&g[16] | &p[38:16]&g[15] | &p[38:15]&g[14] | &p[38:14]&g[13] | &p[38:13]&g[12] | &p[38:12]&g[11] | &p[38:11]&g[10] | &p[38:10]&g[9] | &p[38:9]&g[8] | &p[38:8]&g[7] | &p[38:7]&g[6] | &p[38:6]&g[5] | &p[38:5]&g[4] | &p[38:4]&g[3] | &p[38:3]&g[2] | &p[38:2]&g[1] | &p[38:1]&g[0] | &p[38:0]&c[0];
	assign c[40] = g[39] | &p[39:39]&g[38] | &p[39:38]&g[37] | &p[39:37]&g[36] | &p[39:36]&g[35] | &p[39:35]&g[34] | &p[39:34]&g[33] | &p[39:33]&g[32] | &p[39:32]&g[31] | &p[39:31]&g[30] | &p[39:30]&g[29] | &p[39:29]&g[28] | &p[39:28]&g[27] | &p[39:27]&g[26] | &p[39:26]&g[25] | &p[39:25]&g[24] | &p[39:24]&g[23] | &p[39:23]&g[22] | &p[39:22]&g[21] | &p[39:21]&g[20] | &p[39:20]&g[19] | &p[39:19]&g[18] | &p[39:18]&g[17] | &p[39:17]&g[16] | &p[39:16]&g[15] | &p[39:15]&g[14] | &p[39:14]&g[13] | &p[39:13]&g[12] | &p[39:12]&g[11] | &p[39:11]&g[10] | &p[39:10]&g[9] | &p[39:9]&g[8] | &p[39:8]&g[7] | &p[39:7]&g[6] | &p[39:6]&g[5] | &p[39:5]&g[4] | &p[39:4]&g[3] | &p[39:3]&g[2] | &p[39:2]&g[1] | &p[39:1]&g[0] | &p[39:0]&c[0];
	assign c[41] = g[40] | &p[40:40]&g[39] | &p[40:39]&g[38] | &p[40:38]&g[37] | &p[40:37]&g[36] | &p[40:36]&g[35] | &p[40:35]&g[34] | &p[40:34]&g[33] | &p[40:33]&g[32] | &p[40:32]&g[31] | &p[40:31]&g[30] | &p[40:30]&g[29] | &p[40:29]&g[28] | &p[40:28]&g[27] | &p[40:27]&g[26] | &p[40:26]&g[25] | &p[40:25]&g[24] | &p[40:24]&g[23] | &p[40:23]&g[22] | &p[40:22]&g[21] | &p[40:21]&g[20] | &p[40:20]&g[19] | &p[40:19]&g[18] | &p[40:18]&g[17] | &p[40:17]&g[16] | &p[40:16]&g[15] | &p[40:15]&g[14] | &p[40:14]&g[13] | &p[40:13]&g[12] | &p[40:12]&g[11] | &p[40:11]&g[10] | &p[40:10]&g[9] | &p[40:9]&g[8] | &p[40:8]&g[7] | &p[40:7]&g[6] | &p[40:6]&g[5] | &p[40:5]&g[4] | &p[40:4]&g[3] | &p[40:3]&g[2] | &p[40:2]&g[1] | &p[40:1]&g[0] | &p[40:0]&c[0];
	assign c[42] = g[41] | &p[41:41]&g[40] | &p[41:40]&g[39] | &p[41:39]&g[38] | &p[41:38]&g[37] | &p[41:37]&g[36] | &p[41:36]&g[35] | &p[41:35]&g[34] | &p[41:34]&g[33] | &p[41:33]&g[32] | &p[41:32]&g[31] | &p[41:31]&g[30] | &p[41:30]&g[29] | &p[41:29]&g[28] | &p[41:28]&g[27] | &p[41:27]&g[26] | &p[41:26]&g[25] | &p[41:25]&g[24] | &p[41:24]&g[23] | &p[41:23]&g[22] | &p[41:22]&g[21] | &p[41:21]&g[20] | &p[41:20]&g[19] | &p[41:19]&g[18] | &p[41:18]&g[17] | &p[41:17]&g[16] | &p[41:16]&g[15] | &p[41:15]&g[14] | &p[41:14]&g[13] | &p[41:13]&g[12] | &p[41:12]&g[11] | &p[41:11]&g[10] | &p[41:10]&g[9] | &p[41:9]&g[8] | &p[41:8]&g[7] | &p[41:7]&g[6] | &p[41:6]&g[5] | &p[41:5]&g[4] | &p[41:4]&g[3] | &p[41:3]&g[2] | &p[41:2]&g[1] | &p[41:1]&g[0] | &p[41:0]&c[0];
	assign c[43] = g[42] | &p[42:42]&g[41] | &p[42:41]&g[40] | &p[42:40]&g[39] | &p[42:39]&g[38] | &p[42:38]&g[37] | &p[42:37]&g[36] | &p[42:36]&g[35] | &p[42:35]&g[34] | &p[42:34]&g[33] | &p[42:33]&g[32] | &p[42:32]&g[31] | &p[42:31]&g[30] | &p[42:30]&g[29] | &p[42:29]&g[28] | &p[42:28]&g[27] | &p[42:27]&g[26] | &p[42:26]&g[25] | &p[42:25]&g[24] | &p[42:24]&g[23] | &p[42:23]&g[22] | &p[42:22]&g[21] | &p[42:21]&g[20] | &p[42:20]&g[19] | &p[42:19]&g[18] | &p[42:18]&g[17] | &p[42:17]&g[16] | &p[42:16]&g[15] | &p[42:15]&g[14] | &p[42:14]&g[13] | &p[42:13]&g[12] | &p[42:12]&g[11] | &p[42:11]&g[10] | &p[42:10]&g[9] | &p[42:9]&g[8] | &p[42:8]&g[7] | &p[42:7]&g[6] | &p[42:6]&g[5] | &p[42:5]&g[4] | &p[42:4]&g[3] | &p[42:3]&g[2] | &p[42:2]&g[1] | &p[42:1]&g[0] | &p[42:0]&c[0];
	assign c[44] = g[43] | &p[43:43]&g[42] | &p[43:42]&g[41] | &p[43:41]&g[40] | &p[43:40]&g[39] | &p[43:39]&g[38] | &p[43:38]&g[37] | &p[43:37]&g[36] | &p[43:36]&g[35] | &p[43:35]&g[34] | &p[43:34]&g[33] | &p[43:33]&g[32] | &p[43:32]&g[31] | &p[43:31]&g[30] | &p[43:30]&g[29] | &p[43:29]&g[28] | &p[43:28]&g[27] | &p[43:27]&g[26] | &p[43:26]&g[25] | &p[43:25]&g[24] | &p[43:24]&g[23] | &p[43:23]&g[22] | &p[43:22]&g[21] | &p[43:21]&g[20] | &p[43:20]&g[19] | &p[43:19]&g[18] | &p[43:18]&g[17] | &p[43:17]&g[16] | &p[43:16]&g[15] | &p[43:15]&g[14] | &p[43:14]&g[13] | &p[43:13]&g[12] | &p[43:12]&g[11] | &p[43:11]&g[10] | &p[43:10]&g[9] | &p[43:9]&g[8] | &p[43:8]&g[7] | &p[43:7]&g[6] | &p[43:6]&g[5] | &p[43:5]&g[4] | &p[43:4]&g[3] | &p[43:3]&g[2] | &p[43:2]&g[1] | &p[43:1]&g[0] | &p[43:0]&c[0];
	assign c[45] = g[44] | &p[44:44]&g[43] | &p[44:43]&g[42] | &p[44:42]&g[41] | &p[44:41]&g[40] | &p[44:40]&g[39] | &p[44:39]&g[38] | &p[44:38]&g[37] | &p[44:37]&g[36] | &p[44:36]&g[35] | &p[44:35]&g[34] | &p[44:34]&g[33] | &p[44:33]&g[32] | &p[44:32]&g[31] | &p[44:31]&g[30] | &p[44:30]&g[29] | &p[44:29]&g[28] | &p[44:28]&g[27] | &p[44:27]&g[26] | &p[44:26]&g[25] | &p[44:25]&g[24] | &p[44:24]&g[23] | &p[44:23]&g[22] | &p[44:22]&g[21] | &p[44:21]&g[20] | &p[44:20]&g[19] | &p[44:19]&g[18] | &p[44:18]&g[17] | &p[44:17]&g[16] | &p[44:16]&g[15] | &p[44:15]&g[14] | &p[44:14]&g[13] | &p[44:13]&g[12] | &p[44:12]&g[11] | &p[44:11]&g[10] | &p[44:10]&g[9] | &p[44:9]&g[8] | &p[44:8]&g[7] | &p[44:7]&g[6] | &p[44:6]&g[5] | &p[44:5]&g[4] | &p[44:4]&g[3] | &p[44:3]&g[2] | &p[44:2]&g[1] | &p[44:1]&g[0] | &p[44:0]&c[0];
	assign c[46] = g[45] | &p[45:45]&g[44] | &p[45:44]&g[43] | &p[45:43]&g[42] | &p[45:42]&g[41] | &p[45:41]&g[40] | &p[45:40]&g[39] | &p[45:39]&g[38] | &p[45:38]&g[37] | &p[45:37]&g[36] | &p[45:36]&g[35] | &p[45:35]&g[34] | &p[45:34]&g[33] | &p[45:33]&g[32] | &p[45:32]&g[31] | &p[45:31]&g[30] | &p[45:30]&g[29] | &p[45:29]&g[28] | &p[45:28]&g[27] | &p[45:27]&g[26] | &p[45:26]&g[25] | &p[45:25]&g[24] | &p[45:24]&g[23] | &p[45:23]&g[22] | &p[45:22]&g[21] | &p[45:21]&g[20] | &p[45:20]&g[19] | &p[45:19]&g[18] | &p[45:18]&g[17] | &p[45:17]&g[16] | &p[45:16]&g[15] | &p[45:15]&g[14] | &p[45:14]&g[13] | &p[45:13]&g[12] | &p[45:12]&g[11] | &p[45:11]&g[10] | &p[45:10]&g[9] | &p[45:9]&g[8] | &p[45:8]&g[7] | &p[45:7]&g[6] | &p[45:6]&g[5] | &p[45:5]&g[4] | &p[45:4]&g[3] | &p[45:3]&g[2] | &p[45:2]&g[1] | &p[45:1]&g[0] | &p[45:0]&c[0];
	assign c[47] = g[46] | &p[46:46]&g[45] | &p[46:45]&g[44] | &p[46:44]&g[43] | &p[46:43]&g[42] | &p[46:42]&g[41] | &p[46:41]&g[40] | &p[46:40]&g[39] | &p[46:39]&g[38] | &p[46:38]&g[37] | &p[46:37]&g[36] | &p[46:36]&g[35] | &p[46:35]&g[34] | &p[46:34]&g[33] | &p[46:33]&g[32] | &p[46:32]&g[31] | &p[46:31]&g[30] | &p[46:30]&g[29] | &p[46:29]&g[28] | &p[46:28]&g[27] | &p[46:27]&g[26] | &p[46:26]&g[25] | &p[46:25]&g[24] | &p[46:24]&g[23] | &p[46:23]&g[22] | &p[46:22]&g[21] | &p[46:21]&g[20] | &p[46:20]&g[19] | &p[46:19]&g[18] | &p[46:18]&g[17] | &p[46:17]&g[16] | &p[46:16]&g[15] | &p[46:15]&g[14] | &p[46:14]&g[13] | &p[46:13]&g[12] | &p[46:12]&g[11] | &p[46:11]&g[10] | &p[46:10]&g[9] | &p[46:9]&g[8] | &p[46:8]&g[7] | &p[46:7]&g[6] | &p[46:6]&g[5] | &p[46:5]&g[4] | &p[46:4]&g[3] | &p[46:3]&g[2] | &p[46:2]&g[1] | &p[46:1]&g[0] | &p[46:0]&c[0];
	assign c[48] = g[47] | &p[47:47]&g[46] | &p[47:46]&g[45] | &p[47:45]&g[44] | &p[47:44]&g[43] | &p[47:43]&g[42] | &p[47:42]&g[41] | &p[47:41]&g[40] | &p[47:40]&g[39] | &p[47:39]&g[38] | &p[47:38]&g[37] | &p[47:37]&g[36] | &p[47:36]&g[35] | &p[47:35]&g[34] | &p[47:34]&g[33] | &p[47:33]&g[32] | &p[47:32]&g[31] | &p[47:31]&g[30] | &p[47:30]&g[29] | &p[47:29]&g[28] | &p[47:28]&g[27] | &p[47:27]&g[26] | &p[47:26]&g[25] | &p[47:25]&g[24] | &p[47:24]&g[23] | &p[47:23]&g[22] | &p[47:22]&g[21] | &p[47:21]&g[20] | &p[47:20]&g[19] | &p[47:19]&g[18] | &p[47:18]&g[17] | &p[47:17]&g[16] | &p[47:16]&g[15] | &p[47:15]&g[14] | &p[47:14]&g[13] | &p[47:13]&g[12] | &p[47:12]&g[11] | &p[47:11]&g[10] | &p[47:10]&g[9] | &p[47:9]&g[8] | &p[47:8]&g[7] | &p[47:7]&g[6] | &p[47:6]&g[5] | &p[47:5]&g[4] | &p[47:4]&g[3] | &p[47:3]&g[2] | &p[47:2]&g[1] | &p[47:1]&g[0] | &p[47:0]&c[0];



	assign s = p^c[47:0];

	assign cOut = c[48];

endmodule
