module CLA_64(x, y, cIn, s, cOut);

	input [63:0] x, y;
	input cIn;

	output [63:0] s;
	output cOut;

	wire [63:0] g, p;
	wire [64:0] c;

	assign g = x&y;
	assign p = x^y;

	assign c[0] = cIn;

	assign c[1] = g[0] | &p[0:0]&c[0];
	assign c[2] = g[1] | &p[1:1]&g[0] | &p[1:0]&c[0];
	assign c[3] = g[2] | &p[2:2]&g[1] | &p[2:1]&g[0] | &p[2:0]&c[0];
	assign c[4] = g[3] | &p[3:3]&g[2] | &p[3:2]&g[1] | &p[3:1]&g[0] | &p[3:0]&c[0];
	assign c[5] = g[4] | &p[4:4]&g[3] | &p[4:3]&g[2] | &p[4:2]&g[1] | &p[4:1]&g[0] | &p[4:0]&c[0];
	assign c[6] = g[5] | &p[5:5]&g[4] | &p[5:4]&g[3] | &p[5:3]&g[2] | &p[5:2]&g[1] | &p[5:1]&g[0] | &p[5:0]&c[0];
	assign c[7] = g[6] | &p[6:6]&g[5] | &p[6:5]&g[4] | &p[6:4]&g[3] | &p[6:3]&g[2] | &p[6:2]&g[1] | &p[6:1]&g[0] | &p[6:0]&c[0];
	assign c[8] = g[7] | &p[7:7]&g[6] | &p[7:6]&g[5] | &p[7:5]&g[4] | &p[7:4]&g[3] | &p[7:3]&g[2] | &p[7:2]&g[1] | &p[7:1]&g[0] | &p[7:0]&c[0];
	assign c[9] = g[8] | &p[8:8]&g[7] | &p[8:7]&g[6] | &p[8:6]&g[5] | &p[8:5]&g[4] | &p[8:4]&g[3] | &p[8:3]&g[2] | &p[8:2]&g[1] | &p[8:1]&g[0] | &p[8:0]&c[0];
	assign c[10] = g[9] | &p[9:9]&g[8] | &p[9:8]&g[7] | &p[9:7]&g[6] | &p[9:6]&g[5] | &p[9:5]&g[4] | &p[9:4]&g[3] | &p[9:3]&g[2] | &p[9:2]&g[1] | &p[9:1]&g[0] | &p[9:0]&c[0];
	assign c[11] = g[10] | &p[10:10]&g[9] | &p[10:9]&g[8] | &p[10:8]&g[7] | &p[10:7]&g[6] | &p[10:6]&g[5] | &p[10:5]&g[4] | &p[10:4]&g[3] | &p[10:3]&g[2] | &p[10:2]&g[1] | &p[10:1]&g[0] | &p[10:0]&c[0];
	assign c[12] = g[11] | &p[11:11]&g[10] | &p[11:10]&g[9] | &p[11:9]&g[8] | &p[11:8]&g[7] | &p[11:7]&g[6] | &p[11:6]&g[5] | &p[11:5]&g[4] | &p[11:4]&g[3] | &p[11:3]&g[2] | &p[11:2]&g[1] | &p[11:1]&g[0] | &p[11:0]&c[0];
	assign c[13] = g[12] | &p[12:12]&g[11] | &p[12:11]&g[10] | &p[12:10]&g[9] | &p[12:9]&g[8] | &p[12:8]&g[7] | &p[12:7]&g[6] | &p[12:6]&g[5] | &p[12:5]&g[4] | &p[12:4]&g[3] | &p[12:3]&g[2] | &p[12:2]&g[1] | &p[12:1]&g[0] | &p[12:0]&c[0];
	assign c[14] = g[13] | &p[13:13]&g[12] | &p[13:12]&g[11] | &p[13:11]&g[10] | &p[13:10]&g[9] | &p[13:9]&g[8] | &p[13:8]&g[7] | &p[13:7]&g[6] | &p[13:6]&g[5] | &p[13:5]&g[4] | &p[13:4]&g[3] | &p[13:3]&g[2] | &p[13:2]&g[1] | &p[13:1]&g[0] | &p[13:0]&c[0];
	assign c[15] = g[14] | &p[14:14]&g[13] | &p[14:13]&g[12] | &p[14:12]&g[11] | &p[14:11]&g[10] | &p[14:10]&g[9] | &p[14:9]&g[8] | &p[14:8]&g[7] | &p[14:7]&g[6] | &p[14:6]&g[5] | &p[14:5]&g[4] | &p[14:4]&g[3] | &p[14:3]&g[2] | &p[14:2]&g[1] | &p[14:1]&g[0] | &p[14:0]&c[0];
	assign c[16] = g[15] | &p[15:15]&g[14] | &p[15:14]&g[13] | &p[15:13]&g[12] | &p[15:12]&g[11] | &p[15:11]&g[10] | &p[15:10]&g[9] | &p[15:9]&g[8] | &p[15:8]&g[7] | &p[15:7]&g[6] | &p[15:6]&g[5] | &p[15:5]&g[4] | &p[15:4]&g[3] | &p[15:3]&g[2] | &p[15:2]&g[1] | &p[15:1]&g[0] | &p[15:0]&c[0];
	assign c[17] = g[16] | &p[16:16]&g[15] | &p[16:15]&g[14] | &p[16:14]&g[13] | &p[16:13]&g[12] | &p[16:12]&g[11] | &p[16:11]&g[10] | &p[16:10]&g[9] | &p[16:9]&g[8] | &p[16:8]&g[7] | &p[16:7]&g[6] | &p[16:6]&g[5] | &p[16:5]&g[4] | &p[16:4]&g[3] | &p[16:3]&g[2] | &p[16:2]&g[1] | &p[16:1]&g[0] | &p[16:0]&c[0];
	assign c[18] = g[17] | &p[17:17]&g[16] | &p[17:16]&g[15] | &p[17:15]&g[14] | &p[17:14]&g[13] | &p[17:13]&g[12] | &p[17:12]&g[11] | &p[17:11]&g[10] | &p[17:10]&g[9] | &p[17:9]&g[8] | &p[17:8]&g[7] | &p[17:7]&g[6] | &p[17:6]&g[5] | &p[17:5]&g[4] | &p[17:4]&g[3] | &p[17:3]&g[2] | &p[17:2]&g[1] | &p[17:1]&g[0] | &p[17:0]&c[0];
	assign c[19] = g[18] | &p[18:18]&g[17] | &p[18:17]&g[16] | &p[18:16]&g[15] | &p[18:15]&g[14] | &p[18:14]&g[13] | &p[18:13]&g[12] | &p[18:12]&g[11] | &p[18:11]&g[10] | &p[18:10]&g[9] | &p[18:9]&g[8] | &p[18:8]&g[7] | &p[18:7]&g[6] | &p[18:6]&g[5] | &p[18:5]&g[4] | &p[18:4]&g[3] | &p[18:3]&g[2] | &p[18:2]&g[1] | &p[18:1]&g[0] | &p[18:0]&c[0];
	assign c[20] = g[19] | &p[19:19]&g[18] | &p[19:18]&g[17] | &p[19:17]&g[16] | &p[19:16]&g[15] | &p[19:15]&g[14] | &p[19:14]&g[13] | &p[19:13]&g[12] | &p[19:12]&g[11] | &p[19:11]&g[10] | &p[19:10]&g[9] | &p[19:9]&g[8] | &p[19:8]&g[7] | &p[19:7]&g[6] | &p[19:6]&g[5] | &p[19:5]&g[4] | &p[19:4]&g[3] | &p[19:3]&g[2] | &p[19:2]&g[1] | &p[19:1]&g[0] | &p[19:0]&c[0];
	assign c[21] = g[20] | &p[20:20]&g[19] | &p[20:19]&g[18] | &p[20:18]&g[17] | &p[20:17]&g[16] | &p[20:16]&g[15] | &p[20:15]&g[14] | &p[20:14]&g[13] | &p[20:13]&g[12] | &p[20:12]&g[11] | &p[20:11]&g[10] | &p[20:10]&g[9] | &p[20:9]&g[8] | &p[20:8]&g[7] | &p[20:7]&g[6] | &p[20:6]&g[5] | &p[20:5]&g[4] | &p[20:4]&g[3] | &p[20:3]&g[2] | &p[20:2]&g[1] | &p[20:1]&g[0] | &p[20:0]&c[0];
	assign c[22] = g[21] | &p[21:21]&g[20] | &p[21:20]&g[19] | &p[21:19]&g[18] | &p[21:18]&g[17] | &p[21:17]&g[16] | &p[21:16]&g[15] | &p[21:15]&g[14] | &p[21:14]&g[13] | &p[21:13]&g[12] | &p[21:12]&g[11] | &p[21:11]&g[10] | &p[21:10]&g[9] | &p[21:9]&g[8] | &p[21:8]&g[7] | &p[21:7]&g[6] | &p[21:6]&g[5] | &p[21:5]&g[4] | &p[21:4]&g[3] | &p[21:3]&g[2] | &p[21:2]&g[1] | &p[21:1]&g[0] | &p[21:0]&c[0];
	assign c[23] = g[22] | &p[22:22]&g[21] | &p[22:21]&g[20] | &p[22:20]&g[19] | &p[22:19]&g[18] | &p[22:18]&g[17] | &p[22:17]&g[16] | &p[22:16]&g[15] | &p[22:15]&g[14] | &p[22:14]&g[13] | &p[22:13]&g[12] | &p[22:12]&g[11] | &p[22:11]&g[10] | &p[22:10]&g[9] | &p[22:9]&g[8] | &p[22:8]&g[7] | &p[22:7]&g[6] | &p[22:6]&g[5] | &p[22:5]&g[4] | &p[22:4]&g[3] | &p[22:3]&g[2] | &p[22:2]&g[1] | &p[22:1]&g[0] | &p[22:0]&c[0];
	assign c[24] = g[23] | &p[23:23]&g[22] | &p[23:22]&g[21] | &p[23:21]&g[20] | &p[23:20]&g[19] | &p[23:19]&g[18] | &p[23:18]&g[17] | &p[23:17]&g[16] | &p[23:16]&g[15] | &p[23:15]&g[14] | &p[23:14]&g[13] | &p[23:13]&g[12] | &p[23:12]&g[11] | &p[23:11]&g[10] | &p[23:10]&g[9] | &p[23:9]&g[8] | &p[23:8]&g[7] | &p[23:7]&g[6] | &p[23:6]&g[5] | &p[23:5]&g[4] | &p[23:4]&g[3] | &p[23:3]&g[2] | &p[23:2]&g[1] | &p[23:1]&g[0] | &p[23:0]&c[0];
	assign c[25] = g[24] | &p[24:24]&g[23] | &p[24:23]&g[22] | &p[24:22]&g[21] | &p[24:21]&g[20] | &p[24:20]&g[19] | &p[24:19]&g[18] | &p[24:18]&g[17] | &p[24:17]&g[16] | &p[24:16]&g[15] | &p[24:15]&g[14] | &p[24:14]&g[13] | &p[24:13]&g[12] | &p[24:12]&g[11] | &p[24:11]&g[10] | &p[24:10]&g[9] | &p[24:9]&g[8] | &p[24:8]&g[7] | &p[24:7]&g[6] | &p[24:6]&g[5] | &p[24:5]&g[4] | &p[24:4]&g[3] | &p[24:3]&g[2] | &p[24:2]&g[1] | &p[24:1]&g[0] | &p[24:0]&c[0];
	assign c[26] = g[25] | &p[25:25]&g[24] | &p[25:24]&g[23] | &p[25:23]&g[22] | &p[25:22]&g[21] | &p[25:21]&g[20] | &p[25:20]&g[19] | &p[25:19]&g[18] | &p[25:18]&g[17] | &p[25:17]&g[16] | &p[25:16]&g[15] | &p[25:15]&g[14] | &p[25:14]&g[13] | &p[25:13]&g[12] | &p[25:12]&g[11] | &p[25:11]&g[10] | &p[25:10]&g[9] | &p[25:9]&g[8] | &p[25:8]&g[7] | &p[25:7]&g[6] | &p[25:6]&g[5] | &p[25:5]&g[4] | &p[25:4]&g[3] | &p[25:3]&g[2] | &p[25:2]&g[1] | &p[25:1]&g[0] | &p[25:0]&c[0];
	assign c[27] = g[26] | &p[26:26]&g[25] | &p[26:25]&g[24] | &p[26:24]&g[23] | &p[26:23]&g[22] | &p[26:22]&g[21] | &p[26:21]&g[20] | &p[26:20]&g[19] | &p[26:19]&g[18] | &p[26:18]&g[17] | &p[26:17]&g[16] | &p[26:16]&g[15] | &p[26:15]&g[14] | &p[26:14]&g[13] | &p[26:13]&g[12] | &p[26:12]&g[11] | &p[26:11]&g[10] | &p[26:10]&g[9] | &p[26:9]&g[8] | &p[26:8]&g[7] | &p[26:7]&g[6] | &p[26:6]&g[5] | &p[26:5]&g[4] | &p[26:4]&g[3] | &p[26:3]&g[2] | &p[26:2]&g[1] | &p[26:1]&g[0] | &p[26:0]&c[0];
	assign c[28] = g[27] | &p[27:27]&g[26] | &p[27:26]&g[25] | &p[27:25]&g[24] | &p[27:24]&g[23] | &p[27:23]&g[22] | &p[27:22]&g[21] | &p[27:21]&g[20] | &p[27:20]&g[19] | &p[27:19]&g[18] | &p[27:18]&g[17] | &p[27:17]&g[16] | &p[27:16]&g[15] | &p[27:15]&g[14] | &p[27:14]&g[13] | &p[27:13]&g[12] | &p[27:12]&g[11] | &p[27:11]&g[10] | &p[27:10]&g[9] | &p[27:9]&g[8] | &p[27:8]&g[7] | &p[27:7]&g[6] | &p[27:6]&g[5] | &p[27:5]&g[4] | &p[27:4]&g[3] | &p[27:3]&g[2] | &p[27:2]&g[1] | &p[27:1]&g[0] | &p[27:0]&c[0];
	assign c[29] = g[28] | &p[28:28]&g[27] | &p[28:27]&g[26] | &p[28:26]&g[25] | &p[28:25]&g[24] | &p[28:24]&g[23] | &p[28:23]&g[22] | &p[28:22]&g[21] | &p[28:21]&g[20] | &p[28:20]&g[19] | &p[28:19]&g[18] | &p[28:18]&g[17] | &p[28:17]&g[16] | &p[28:16]&g[15] | &p[28:15]&g[14] | &p[28:14]&g[13] | &p[28:13]&g[12] | &p[28:12]&g[11] | &p[28:11]&g[10] | &p[28:10]&g[9] | &p[28:9]&g[8] | &p[28:8]&g[7] | &p[28:7]&g[6] | &p[28:6]&g[5] | &p[28:5]&g[4] | &p[28:4]&g[3] | &p[28:3]&g[2] | &p[28:2]&g[1] | &p[28:1]&g[0] | &p[28:0]&c[0];
	assign c[30] = g[29] | &p[29:29]&g[28] | &p[29:28]&g[27] | &p[29:27]&g[26] | &p[29:26]&g[25] | &p[29:25]&g[24] | &p[29:24]&g[23] | &p[29:23]&g[22] | &p[29:22]&g[21] | &p[29:21]&g[20] | &p[29:20]&g[19] | &p[29:19]&g[18] | &p[29:18]&g[17] | &p[29:17]&g[16] | &p[29:16]&g[15] | &p[29:15]&g[14] | &p[29:14]&g[13] | &p[29:13]&g[12] | &p[29:12]&g[11] | &p[29:11]&g[10] | &p[29:10]&g[9] | &p[29:9]&g[8] | &p[29:8]&g[7] | &p[29:7]&g[6] | &p[29:6]&g[5] | &p[29:5]&g[4] | &p[29:4]&g[3] | &p[29:3]&g[2] | &p[29:2]&g[1] | &p[29:1]&g[0] | &p[29:0]&c[0];
	assign c[31] = g[30] | &p[30:30]&g[29] | &p[30:29]&g[28] | &p[30:28]&g[27] | &p[30:27]&g[26] | &p[30:26]&g[25] | &p[30:25]&g[24] | &p[30:24]&g[23] | &p[30:23]&g[22] | &p[30:22]&g[21] | &p[30:21]&g[20] | &p[30:20]&g[19] | &p[30:19]&g[18] | &p[30:18]&g[17] | &p[30:17]&g[16] | &p[30:16]&g[15] | &p[30:15]&g[14] | &p[30:14]&g[13] | &p[30:13]&g[12] | &p[30:12]&g[11] | &p[30:11]&g[10] | &p[30:10]&g[9] | &p[30:9]&g[8] | &p[30:8]&g[7] | &p[30:7]&g[6] | &p[30:6]&g[5] | &p[30:5]&g[4] | &p[30:4]&g[3] | &p[30:3]&g[2] | &p[30:2]&g[1] | &p[30:1]&g[0] | &p[30:0]&c[0];
	assign c[32] = g[31] | &p[31:31]&g[30] | &p[31:30]&g[29] | &p[31:29]&g[28] | &p[31:28]&g[27] | &p[31:27]&g[26] | &p[31:26]&g[25] | &p[31:25]&g[24] | &p[31:24]&g[23] | &p[31:23]&g[22] | &p[31:22]&g[21] | &p[31:21]&g[20] | &p[31:20]&g[19] | &p[31:19]&g[18] | &p[31:18]&g[17] | &p[31:17]&g[16] | &p[31:16]&g[15] | &p[31:15]&g[14] | &p[31:14]&g[13] | &p[31:13]&g[12] | &p[31:12]&g[11] | &p[31:11]&g[10] | &p[31:10]&g[9] | &p[31:9]&g[8] | &p[31:8]&g[7] | &p[31:7]&g[6] | &p[31:6]&g[5] | &p[31:5]&g[4] | &p[31:4]&g[3] | &p[31:3]&g[2] | &p[31:2]&g[1] | &p[31:1]&g[0] | &p[31:0]&c[0];
	assign c[33] = g[32] | &p[32:32]&g[31] | &p[32:31]&g[30] | &p[32:30]&g[29] | &p[32:29]&g[28] | &p[32:28]&g[27] | &p[32:27]&g[26] | &p[32:26]&g[25] | &p[32:25]&g[24] | &p[32:24]&g[23] | &p[32:23]&g[22] | &p[32:22]&g[21] | &p[32:21]&g[20] | &p[32:20]&g[19] | &p[32:19]&g[18] | &p[32:18]&g[17] | &p[32:17]&g[16] | &p[32:16]&g[15] | &p[32:15]&g[14] | &p[32:14]&g[13] | &p[32:13]&g[12] | &p[32:12]&g[11] | &p[32:11]&g[10] | &p[32:10]&g[9] | &p[32:9]&g[8] | &p[32:8]&g[7] | &p[32:7]&g[6] | &p[32:6]&g[5] | &p[32:5]&g[4] | &p[32:4]&g[3] | &p[32:3]&g[2] | &p[32:2]&g[1] | &p[32:1]&g[0] | &p[32:0]&c[0];
	assign c[34] = g[33] | &p[33:33]&g[32] | &p[33:32]&g[31] | &p[33:31]&g[30] | &p[33:30]&g[29] | &p[33:29]&g[28] | &p[33:28]&g[27] | &p[33:27]&g[26] | &p[33:26]&g[25] | &p[33:25]&g[24] | &p[33:24]&g[23] | &p[33:23]&g[22] | &p[33:22]&g[21] | &p[33:21]&g[20] | &p[33:20]&g[19] | &p[33:19]&g[18] | &p[33:18]&g[17] | &p[33:17]&g[16] | &p[33:16]&g[15] | &p[33:15]&g[14] | &p[33:14]&g[13] | &p[33:13]&g[12] | &p[33:12]&g[11] | &p[33:11]&g[10] | &p[33:10]&g[9] | &p[33:9]&g[8] | &p[33:8]&g[7] | &p[33:7]&g[6] | &p[33:6]&g[5] | &p[33:5]&g[4] | &p[33:4]&g[3] | &p[33:3]&g[2] | &p[33:2]&g[1] | &p[33:1]&g[0] | &p[33:0]&c[0];
	assign c[35] = g[34] | &p[34:34]&g[33] | &p[34:33]&g[32] | &p[34:32]&g[31] | &p[34:31]&g[30] | &p[34:30]&g[29] | &p[34:29]&g[28] | &p[34:28]&g[27] | &p[34:27]&g[26] | &p[34:26]&g[25] | &p[34:25]&g[24] | &p[34:24]&g[23] | &p[34:23]&g[22] | &p[34:22]&g[21] | &p[34:21]&g[20] | &p[34:20]&g[19] | &p[34:19]&g[18] | &p[34:18]&g[17] | &p[34:17]&g[16] | &p[34:16]&g[15] | &p[34:15]&g[14] | &p[34:14]&g[13] | &p[34:13]&g[12] | &p[34:12]&g[11] | &p[34:11]&g[10] | &p[34:10]&g[9] | &p[34:9]&g[8] | &p[34:8]&g[7] | &p[34:7]&g[6] | &p[34:6]&g[5] | &p[34:5]&g[4] | &p[34:4]&g[3] | &p[34:3]&g[2] | &p[34:2]&g[1] | &p[34:1]&g[0] | &p[34:0]&c[0];
	assign c[36] = g[35] | &p[35:35]&g[34] | &p[35:34]&g[33] | &p[35:33]&g[32] | &p[35:32]&g[31] | &p[35:31]&g[30] | &p[35:30]&g[29] | &p[35:29]&g[28] | &p[35:28]&g[27] | &p[35:27]&g[26] | &p[35:26]&g[25] | &p[35:25]&g[24] | &p[35:24]&g[23] | &p[35:23]&g[22] | &p[35:22]&g[21] | &p[35:21]&g[20] | &p[35:20]&g[19] | &p[35:19]&g[18] | &p[35:18]&g[17] | &p[35:17]&g[16] | &p[35:16]&g[15] | &p[35:15]&g[14] | &p[35:14]&g[13] | &p[35:13]&g[12] | &p[35:12]&g[11] | &p[35:11]&g[10] | &p[35:10]&g[9] | &p[35:9]&g[8] | &p[35:8]&g[7] | &p[35:7]&g[6] | &p[35:6]&g[5] | &p[35:5]&g[4] | &p[35:4]&g[3] | &p[35:3]&g[2] | &p[35:2]&g[1] | &p[35:1]&g[0] | &p[35:0]&c[0];
	assign c[37] = g[36] | &p[36:36]&g[35] | &p[36:35]&g[34] | &p[36:34]&g[33] | &p[36:33]&g[32] | &p[36:32]&g[31] | &p[36:31]&g[30] | &p[36:30]&g[29] | &p[36:29]&g[28] | &p[36:28]&g[27] | &p[36:27]&g[26] | &p[36:26]&g[25] | &p[36:25]&g[24] | &p[36:24]&g[23] | &p[36:23]&g[22] | &p[36:22]&g[21] | &p[36:21]&g[20] | &p[36:20]&g[19] | &p[36:19]&g[18] | &p[36:18]&g[17] | &p[36:17]&g[16] | &p[36:16]&g[15] | &p[36:15]&g[14] | &p[36:14]&g[13] | &p[36:13]&g[12] | &p[36:12]&g[11] | &p[36:11]&g[10] | &p[36:10]&g[9] | &p[36:9]&g[8] | &p[36:8]&g[7] | &p[36:7]&g[6] | &p[36:6]&g[5] | &p[36:5]&g[4] | &p[36:4]&g[3] | &p[36:3]&g[2] | &p[36:2]&g[1] | &p[36:1]&g[0] | &p[36:0]&c[0];
	assign c[38] = g[37] | &p[37:37]&g[36] | &p[37:36]&g[35] | &p[37:35]&g[34] | &p[37:34]&g[33] | &p[37:33]&g[32] | &p[37:32]&g[31] | &p[37:31]&g[30] | &p[37:30]&g[29] | &p[37:29]&g[28] | &p[37:28]&g[27] | &p[37:27]&g[26] | &p[37:26]&g[25] | &p[37:25]&g[24] | &p[37:24]&g[23] | &p[37:23]&g[22] | &p[37:22]&g[21] | &p[37:21]&g[20] | &p[37:20]&g[19] | &p[37:19]&g[18] | &p[37:18]&g[17] | &p[37:17]&g[16] | &p[37:16]&g[15] | &p[37:15]&g[14] | &p[37:14]&g[13] | &p[37:13]&g[12] | &p[37:12]&g[11] | &p[37:11]&g[10] | &p[37:10]&g[9] | &p[37:9]&g[8] | &p[37:8]&g[7] | &p[37:7]&g[6] | &p[37:6]&g[5] | &p[37:5]&g[4] | &p[37:4]&g[3] | &p[37:3]&g[2] | &p[37:2]&g[1] | &p[37:1]&g[0] | &p[37:0]&c[0];
	assign c[39] = g[38] | &p[38:38]&g[37] | &p[38:37]&g[36] | &p[38:36]&g[35] | &p[38:35]&g[34] | &p[38:34]&g[33] | &p[38:33]&g[32] | &p[38:32]&g[31] | &p[38:31]&g[30] | &p[38:30]&g[29] | &p[38:29]&g[28] | &p[38:28]&g[27] | &p[38:27]&g[26] | &p[38:26]&g[25] | &p[38:25]&g[24] | &p[38:24]&g[23] | &p[38:23]&g[22] | &p[38:22]&g[21] | &p[38:21]&g[20] | &p[38:20]&g[19] | &p[38:19]&g[18] | &p[38:18]&g[17] | &p[38:17]&g[16] | &p[38:16]&g[15] | &p[38:15]&g[14] | &p[38:14]&g[13] | &p[38:13]&g[12] | &p[38:12]&g[11] | &p[38:11]&g[10] | &p[38:10]&g[9] | &p[38:9]&g[8] | &p[38:8]&g[7] | &p[38:7]&g[6] | &p[38:6]&g[5] | &p[38:5]&g[4] | &p[38:4]&g[3] | &p[38:3]&g[2] | &p[38:2]&g[1] | &p[38:1]&g[0] | &p[38:0]&c[0];
	assign c[40] = g[39] | &p[39:39]&g[38] | &p[39:38]&g[37] | &p[39:37]&g[36] | &p[39:36]&g[35] | &p[39:35]&g[34] | &p[39:34]&g[33] | &p[39:33]&g[32] | &p[39:32]&g[31] | &p[39:31]&g[30] | &p[39:30]&g[29] | &p[39:29]&g[28] | &p[39:28]&g[27] | &p[39:27]&g[26] | &p[39:26]&g[25] | &p[39:25]&g[24] | &p[39:24]&g[23] | &p[39:23]&g[22] | &p[39:22]&g[21] | &p[39:21]&g[20] | &p[39:20]&g[19] | &p[39:19]&g[18] | &p[39:18]&g[17] | &p[39:17]&g[16] | &p[39:16]&g[15] | &p[39:15]&g[14] | &p[39:14]&g[13] | &p[39:13]&g[12] | &p[39:12]&g[11] | &p[39:11]&g[10] | &p[39:10]&g[9] | &p[39:9]&g[8] | &p[39:8]&g[7] | &p[39:7]&g[6] | &p[39:6]&g[5] | &p[39:5]&g[4] | &p[39:4]&g[3] | &p[39:3]&g[2] | &p[39:2]&g[1] | &p[39:1]&g[0] | &p[39:0]&c[0];
	assign c[41] = g[40] | &p[40:40]&g[39] | &p[40:39]&g[38] | &p[40:38]&g[37] | &p[40:37]&g[36] | &p[40:36]&g[35] | &p[40:35]&g[34] | &p[40:34]&g[33] | &p[40:33]&g[32] | &p[40:32]&g[31] | &p[40:31]&g[30] | &p[40:30]&g[29] | &p[40:29]&g[28] | &p[40:28]&g[27] | &p[40:27]&g[26] | &p[40:26]&g[25] | &p[40:25]&g[24] | &p[40:24]&g[23] | &p[40:23]&g[22] | &p[40:22]&g[21] | &p[40:21]&g[20] | &p[40:20]&g[19] | &p[40:19]&g[18] | &p[40:18]&g[17] | &p[40:17]&g[16] | &p[40:16]&g[15] | &p[40:15]&g[14] | &p[40:14]&g[13] | &p[40:13]&g[12] | &p[40:12]&g[11] | &p[40:11]&g[10] | &p[40:10]&g[9] | &p[40:9]&g[8] | &p[40:8]&g[7] | &p[40:7]&g[6] | &p[40:6]&g[5] | &p[40:5]&g[4] | &p[40:4]&g[3] | &p[40:3]&g[2] | &p[40:2]&g[1] | &p[40:1]&g[0] | &p[40:0]&c[0];
	assign c[42] = g[41] | &p[41:41]&g[40] | &p[41:40]&g[39] | &p[41:39]&g[38] | &p[41:38]&g[37] | &p[41:37]&g[36] | &p[41:36]&g[35] | &p[41:35]&g[34] | &p[41:34]&g[33] | &p[41:33]&g[32] | &p[41:32]&g[31] | &p[41:31]&g[30] | &p[41:30]&g[29] | &p[41:29]&g[28] | &p[41:28]&g[27] | &p[41:27]&g[26] | &p[41:26]&g[25] | &p[41:25]&g[24] | &p[41:24]&g[23] | &p[41:23]&g[22] | &p[41:22]&g[21] | &p[41:21]&g[20] | &p[41:20]&g[19] | &p[41:19]&g[18] | &p[41:18]&g[17] | &p[41:17]&g[16] | &p[41:16]&g[15] | &p[41:15]&g[14] | &p[41:14]&g[13] | &p[41:13]&g[12] | &p[41:12]&g[11] | &p[41:11]&g[10] | &p[41:10]&g[9] | &p[41:9]&g[8] | &p[41:8]&g[7] | &p[41:7]&g[6] | &p[41:6]&g[5] | &p[41:5]&g[4] | &p[41:4]&g[3] | &p[41:3]&g[2] | &p[41:2]&g[1] | &p[41:1]&g[0] | &p[41:0]&c[0];
	assign c[43] = g[42] | &p[42:42]&g[41] | &p[42:41]&g[40] | &p[42:40]&g[39] | &p[42:39]&g[38] | &p[42:38]&g[37] | &p[42:37]&g[36] | &p[42:36]&g[35] | &p[42:35]&g[34] | &p[42:34]&g[33] | &p[42:33]&g[32] | &p[42:32]&g[31] | &p[42:31]&g[30] | &p[42:30]&g[29] | &p[42:29]&g[28] | &p[42:28]&g[27] | &p[42:27]&g[26] | &p[42:26]&g[25] | &p[42:25]&g[24] | &p[42:24]&g[23] | &p[42:23]&g[22] | &p[42:22]&g[21] | &p[42:21]&g[20] | &p[42:20]&g[19] | &p[42:19]&g[18] | &p[42:18]&g[17] | &p[42:17]&g[16] | &p[42:16]&g[15] | &p[42:15]&g[14] | &p[42:14]&g[13] | &p[42:13]&g[12] | &p[42:12]&g[11] | &p[42:11]&g[10] | &p[42:10]&g[9] | &p[42:9]&g[8] | &p[42:8]&g[7] | &p[42:7]&g[6] | &p[42:6]&g[5] | &p[42:5]&g[4] | &p[42:4]&g[3] | &p[42:3]&g[2] | &p[42:2]&g[1] | &p[42:1]&g[0] | &p[42:0]&c[0];
	assign c[44] = g[43] | &p[43:43]&g[42] | &p[43:42]&g[41] | &p[43:41]&g[40] | &p[43:40]&g[39] | &p[43:39]&g[38] | &p[43:38]&g[37] | &p[43:37]&g[36] | &p[43:36]&g[35] | &p[43:35]&g[34] | &p[43:34]&g[33] | &p[43:33]&g[32] | &p[43:32]&g[31] | &p[43:31]&g[30] | &p[43:30]&g[29] | &p[43:29]&g[28] | &p[43:28]&g[27] | &p[43:27]&g[26] | &p[43:26]&g[25] | &p[43:25]&g[24] | &p[43:24]&g[23] | &p[43:23]&g[22] | &p[43:22]&g[21] | &p[43:21]&g[20] | &p[43:20]&g[19] | &p[43:19]&g[18] | &p[43:18]&g[17] | &p[43:17]&g[16] | &p[43:16]&g[15] | &p[43:15]&g[14] | &p[43:14]&g[13] | &p[43:13]&g[12] | &p[43:12]&g[11] | &p[43:11]&g[10] | &p[43:10]&g[9] | &p[43:9]&g[8] | &p[43:8]&g[7] | &p[43:7]&g[6] | &p[43:6]&g[5] | &p[43:5]&g[4] | &p[43:4]&g[3] | &p[43:3]&g[2] | &p[43:2]&g[1] | &p[43:1]&g[0] | &p[43:0]&c[0];
	assign c[45] = g[44] | &p[44:44]&g[43] | &p[44:43]&g[42] | &p[44:42]&g[41] | &p[44:41]&g[40] | &p[44:40]&g[39] | &p[44:39]&g[38] | &p[44:38]&g[37] | &p[44:37]&g[36] | &p[44:36]&g[35] | &p[44:35]&g[34] | &p[44:34]&g[33] | &p[44:33]&g[32] | &p[44:32]&g[31] | &p[44:31]&g[30] | &p[44:30]&g[29] | &p[44:29]&g[28] | &p[44:28]&g[27] | &p[44:27]&g[26] | &p[44:26]&g[25] | &p[44:25]&g[24] | &p[44:24]&g[23] | &p[44:23]&g[22] | &p[44:22]&g[21] | &p[44:21]&g[20] | &p[44:20]&g[19] | &p[44:19]&g[18] | &p[44:18]&g[17] | &p[44:17]&g[16] | &p[44:16]&g[15] | &p[44:15]&g[14] | &p[44:14]&g[13] | &p[44:13]&g[12] | &p[44:12]&g[11] | &p[44:11]&g[10] | &p[44:10]&g[9] | &p[44:9]&g[8] | &p[44:8]&g[7] | &p[44:7]&g[6] | &p[44:6]&g[5] | &p[44:5]&g[4] | &p[44:4]&g[3] | &p[44:3]&g[2] | &p[44:2]&g[1] | &p[44:1]&g[0] | &p[44:0]&c[0];
	assign c[46] = g[45] | &p[45:45]&g[44] | &p[45:44]&g[43] | &p[45:43]&g[42] | &p[45:42]&g[41] | &p[45:41]&g[40] | &p[45:40]&g[39] | &p[45:39]&g[38] | &p[45:38]&g[37] | &p[45:37]&g[36] | &p[45:36]&g[35] | &p[45:35]&g[34] | &p[45:34]&g[33] | &p[45:33]&g[32] | &p[45:32]&g[31] | &p[45:31]&g[30] | &p[45:30]&g[29] | &p[45:29]&g[28] | &p[45:28]&g[27] | &p[45:27]&g[26] | &p[45:26]&g[25] | &p[45:25]&g[24] | &p[45:24]&g[23] | &p[45:23]&g[22] | &p[45:22]&g[21] | &p[45:21]&g[20] | &p[45:20]&g[19] | &p[45:19]&g[18] | &p[45:18]&g[17] | &p[45:17]&g[16] | &p[45:16]&g[15] | &p[45:15]&g[14] | &p[45:14]&g[13] | &p[45:13]&g[12] | &p[45:12]&g[11] | &p[45:11]&g[10] | &p[45:10]&g[9] | &p[45:9]&g[8] | &p[45:8]&g[7] | &p[45:7]&g[6] | &p[45:6]&g[5] | &p[45:5]&g[4] | &p[45:4]&g[3] | &p[45:3]&g[2] | &p[45:2]&g[1] | &p[45:1]&g[0] | &p[45:0]&c[0];
	assign c[47] = g[46] | &p[46:46]&g[45] | &p[46:45]&g[44] | &p[46:44]&g[43] | &p[46:43]&g[42] | &p[46:42]&g[41] | &p[46:41]&g[40] | &p[46:40]&g[39] | &p[46:39]&g[38] | &p[46:38]&g[37] | &p[46:37]&g[36] | &p[46:36]&g[35] | &p[46:35]&g[34] | &p[46:34]&g[33] | &p[46:33]&g[32] | &p[46:32]&g[31] | &p[46:31]&g[30] | &p[46:30]&g[29] | &p[46:29]&g[28] | &p[46:28]&g[27] | &p[46:27]&g[26] | &p[46:26]&g[25] | &p[46:25]&g[24] | &p[46:24]&g[23] | &p[46:23]&g[22] | &p[46:22]&g[21] | &p[46:21]&g[20] | &p[46:20]&g[19] | &p[46:19]&g[18] | &p[46:18]&g[17] | &p[46:17]&g[16] | &p[46:16]&g[15] | &p[46:15]&g[14] | &p[46:14]&g[13] | &p[46:13]&g[12] | &p[46:12]&g[11] | &p[46:11]&g[10] | &p[46:10]&g[9] | &p[46:9]&g[8] | &p[46:8]&g[7] | &p[46:7]&g[6] | &p[46:6]&g[5] | &p[46:5]&g[4] | &p[46:4]&g[3] | &p[46:3]&g[2] | &p[46:2]&g[1] | &p[46:1]&g[0] | &p[46:0]&c[0];
	assign c[48] = g[47] | &p[47:47]&g[46] | &p[47:46]&g[45] | &p[47:45]&g[44] | &p[47:44]&g[43] | &p[47:43]&g[42] | &p[47:42]&g[41] | &p[47:41]&g[40] | &p[47:40]&g[39] | &p[47:39]&g[38] | &p[47:38]&g[37] | &p[47:37]&g[36] | &p[47:36]&g[35] | &p[47:35]&g[34] | &p[47:34]&g[33] | &p[47:33]&g[32] | &p[47:32]&g[31] | &p[47:31]&g[30] | &p[47:30]&g[29] | &p[47:29]&g[28] | &p[47:28]&g[27] | &p[47:27]&g[26] | &p[47:26]&g[25] | &p[47:25]&g[24] | &p[47:24]&g[23] | &p[47:23]&g[22] | &p[47:22]&g[21] | &p[47:21]&g[20] | &p[47:20]&g[19] | &p[47:19]&g[18] | &p[47:18]&g[17] | &p[47:17]&g[16] | &p[47:16]&g[15] | &p[47:15]&g[14] | &p[47:14]&g[13] | &p[47:13]&g[12] | &p[47:12]&g[11] | &p[47:11]&g[10] | &p[47:10]&g[9] | &p[47:9]&g[8] | &p[47:8]&g[7] | &p[47:7]&g[6] | &p[47:6]&g[5] | &p[47:5]&g[4] | &p[47:4]&g[3] | &p[47:3]&g[2] | &p[47:2]&g[1] | &p[47:1]&g[0] | &p[47:0]&c[0];
	assign c[49] = g[48] | &p[48:48]&g[47] | &p[48:47]&g[46] | &p[48:46]&g[45] | &p[48:45]&g[44] | &p[48:44]&g[43] | &p[48:43]&g[42] | &p[48:42]&g[41] | &p[48:41]&g[40] | &p[48:40]&g[39] | &p[48:39]&g[38] | &p[48:38]&g[37] | &p[48:37]&g[36] | &p[48:36]&g[35] | &p[48:35]&g[34] | &p[48:34]&g[33] | &p[48:33]&g[32] | &p[48:32]&g[31] | &p[48:31]&g[30] | &p[48:30]&g[29] | &p[48:29]&g[28] | &p[48:28]&g[27] | &p[48:27]&g[26] | &p[48:26]&g[25] | &p[48:25]&g[24] | &p[48:24]&g[23] | &p[48:23]&g[22] | &p[48:22]&g[21] | &p[48:21]&g[20] | &p[48:20]&g[19] | &p[48:19]&g[18] | &p[48:18]&g[17] | &p[48:17]&g[16] | &p[48:16]&g[15] | &p[48:15]&g[14] | &p[48:14]&g[13] | &p[48:13]&g[12] | &p[48:12]&g[11] | &p[48:11]&g[10] | &p[48:10]&g[9] | &p[48:9]&g[8] | &p[48:8]&g[7] | &p[48:7]&g[6] | &p[48:6]&g[5] | &p[48:5]&g[4] | &p[48:4]&g[3] | &p[48:3]&g[2] | &p[48:2]&g[1] | &p[48:1]&g[0] | &p[48:0]&c[0];
	assign c[50] = g[49] | &p[49:49]&g[48] | &p[49:48]&g[47] | &p[49:47]&g[46] | &p[49:46]&g[45] | &p[49:45]&g[44] | &p[49:44]&g[43] | &p[49:43]&g[42] | &p[49:42]&g[41] | &p[49:41]&g[40] | &p[49:40]&g[39] | &p[49:39]&g[38] | &p[49:38]&g[37] | &p[49:37]&g[36] | &p[49:36]&g[35] | &p[49:35]&g[34] | &p[49:34]&g[33] | &p[49:33]&g[32] | &p[49:32]&g[31] | &p[49:31]&g[30] | &p[49:30]&g[29] | &p[49:29]&g[28] | &p[49:28]&g[27] | &p[49:27]&g[26] | &p[49:26]&g[25] | &p[49:25]&g[24] | &p[49:24]&g[23] | &p[49:23]&g[22] | &p[49:22]&g[21] | &p[49:21]&g[20] | &p[49:20]&g[19] | &p[49:19]&g[18] | &p[49:18]&g[17] | &p[49:17]&g[16] | &p[49:16]&g[15] | &p[49:15]&g[14] | &p[49:14]&g[13] | &p[49:13]&g[12] | &p[49:12]&g[11] | &p[49:11]&g[10] | &p[49:10]&g[9] | &p[49:9]&g[8] | &p[49:8]&g[7] | &p[49:7]&g[6] | &p[49:6]&g[5] | &p[49:5]&g[4] | &p[49:4]&g[3] | &p[49:3]&g[2] | &p[49:2]&g[1] | &p[49:1]&g[0] | &p[49:0]&c[0];
	assign c[51] = g[50] | &p[50:50]&g[49] | &p[50:49]&g[48] | &p[50:48]&g[47] | &p[50:47]&g[46] | &p[50:46]&g[45] | &p[50:45]&g[44] | &p[50:44]&g[43] | &p[50:43]&g[42] | &p[50:42]&g[41] | &p[50:41]&g[40] | &p[50:40]&g[39] | &p[50:39]&g[38] | &p[50:38]&g[37] | &p[50:37]&g[36] | &p[50:36]&g[35] | &p[50:35]&g[34] | &p[50:34]&g[33] | &p[50:33]&g[32] | &p[50:32]&g[31] | &p[50:31]&g[30] | &p[50:30]&g[29] | &p[50:29]&g[28] | &p[50:28]&g[27] | &p[50:27]&g[26] | &p[50:26]&g[25] | &p[50:25]&g[24] | &p[50:24]&g[23] | &p[50:23]&g[22] | &p[50:22]&g[21] | &p[50:21]&g[20] | &p[50:20]&g[19] | &p[50:19]&g[18] | &p[50:18]&g[17] | &p[50:17]&g[16] | &p[50:16]&g[15] | &p[50:15]&g[14] | &p[50:14]&g[13] | &p[50:13]&g[12] | &p[50:12]&g[11] | &p[50:11]&g[10] | &p[50:10]&g[9] | &p[50:9]&g[8] | &p[50:8]&g[7] | &p[50:7]&g[6] | &p[50:6]&g[5] | &p[50:5]&g[4] | &p[50:4]&g[3] | &p[50:3]&g[2] | &p[50:2]&g[1] | &p[50:1]&g[0] | &p[50:0]&c[0];
	assign c[52] = g[51] | &p[51:51]&g[50] | &p[51:50]&g[49] | &p[51:49]&g[48] | &p[51:48]&g[47] | &p[51:47]&g[46] | &p[51:46]&g[45] | &p[51:45]&g[44] | &p[51:44]&g[43] | &p[51:43]&g[42] | &p[51:42]&g[41] | &p[51:41]&g[40] | &p[51:40]&g[39] | &p[51:39]&g[38] | &p[51:38]&g[37] | &p[51:37]&g[36] | &p[51:36]&g[35] | &p[51:35]&g[34] | &p[51:34]&g[33] | &p[51:33]&g[32] | &p[51:32]&g[31] | &p[51:31]&g[30] | &p[51:30]&g[29] | &p[51:29]&g[28] | &p[51:28]&g[27] | &p[51:27]&g[26] | &p[51:26]&g[25] | &p[51:25]&g[24] | &p[51:24]&g[23] | &p[51:23]&g[22] | &p[51:22]&g[21] | &p[51:21]&g[20] | &p[51:20]&g[19] | &p[51:19]&g[18] | &p[51:18]&g[17] | &p[51:17]&g[16] | &p[51:16]&g[15] | &p[51:15]&g[14] | &p[51:14]&g[13] | &p[51:13]&g[12] | &p[51:12]&g[11] | &p[51:11]&g[10] | &p[51:10]&g[9] | &p[51:9]&g[8] | &p[51:8]&g[7] | &p[51:7]&g[6] | &p[51:6]&g[5] | &p[51:5]&g[4] | &p[51:4]&g[3] | &p[51:3]&g[2] | &p[51:2]&g[1] | &p[51:1]&g[0] | &p[51:0]&c[0];
	assign c[53] = g[52] | &p[52:52]&g[51] | &p[52:51]&g[50] | &p[52:50]&g[49] | &p[52:49]&g[48] | &p[52:48]&g[47] | &p[52:47]&g[46] | &p[52:46]&g[45] | &p[52:45]&g[44] | &p[52:44]&g[43] | &p[52:43]&g[42] | &p[52:42]&g[41] | &p[52:41]&g[40] | &p[52:40]&g[39] | &p[52:39]&g[38] | &p[52:38]&g[37] | &p[52:37]&g[36] | &p[52:36]&g[35] | &p[52:35]&g[34] | &p[52:34]&g[33] | &p[52:33]&g[32] | &p[52:32]&g[31] | &p[52:31]&g[30] | &p[52:30]&g[29] | &p[52:29]&g[28] | &p[52:28]&g[27] | &p[52:27]&g[26] | &p[52:26]&g[25] | &p[52:25]&g[24] | &p[52:24]&g[23] | &p[52:23]&g[22] | &p[52:22]&g[21] | &p[52:21]&g[20] | &p[52:20]&g[19] | &p[52:19]&g[18] | &p[52:18]&g[17] | &p[52:17]&g[16] | &p[52:16]&g[15] | &p[52:15]&g[14] | &p[52:14]&g[13] | &p[52:13]&g[12] | &p[52:12]&g[11] | &p[52:11]&g[10] | &p[52:10]&g[9] | &p[52:9]&g[8] | &p[52:8]&g[7] | &p[52:7]&g[6] | &p[52:6]&g[5] | &p[52:5]&g[4] | &p[52:4]&g[3] | &p[52:3]&g[2] | &p[52:2]&g[1] | &p[52:1]&g[0] | &p[52:0]&c[0];
	assign c[54] = g[53] | &p[53:53]&g[52] | &p[53:52]&g[51] | &p[53:51]&g[50] | &p[53:50]&g[49] | &p[53:49]&g[48] | &p[53:48]&g[47] | &p[53:47]&g[46] | &p[53:46]&g[45] | &p[53:45]&g[44] | &p[53:44]&g[43] | &p[53:43]&g[42] | &p[53:42]&g[41] | &p[53:41]&g[40] | &p[53:40]&g[39] | &p[53:39]&g[38] | &p[53:38]&g[37] | &p[53:37]&g[36] | &p[53:36]&g[35] | &p[53:35]&g[34] | &p[53:34]&g[33] | &p[53:33]&g[32] | &p[53:32]&g[31] | &p[53:31]&g[30] | &p[53:30]&g[29] | &p[53:29]&g[28] | &p[53:28]&g[27] | &p[53:27]&g[26] | &p[53:26]&g[25] | &p[53:25]&g[24] | &p[53:24]&g[23] | &p[53:23]&g[22] | &p[53:22]&g[21] | &p[53:21]&g[20] | &p[53:20]&g[19] | &p[53:19]&g[18] | &p[53:18]&g[17] | &p[53:17]&g[16] | &p[53:16]&g[15] | &p[53:15]&g[14] | &p[53:14]&g[13] | &p[53:13]&g[12] | &p[53:12]&g[11] | &p[53:11]&g[10] | &p[53:10]&g[9] | &p[53:9]&g[8] | &p[53:8]&g[7] | &p[53:7]&g[6] | &p[53:6]&g[5] | &p[53:5]&g[4] | &p[53:4]&g[3] | &p[53:3]&g[2] | &p[53:2]&g[1] | &p[53:1]&g[0] | &p[53:0]&c[0];
	assign c[55] = g[54] | &p[54:54]&g[53] | &p[54:53]&g[52] | &p[54:52]&g[51] | &p[54:51]&g[50] | &p[54:50]&g[49] | &p[54:49]&g[48] | &p[54:48]&g[47] | &p[54:47]&g[46] | &p[54:46]&g[45] | &p[54:45]&g[44] | &p[54:44]&g[43] | &p[54:43]&g[42] | &p[54:42]&g[41] | &p[54:41]&g[40] | &p[54:40]&g[39] | &p[54:39]&g[38] | &p[54:38]&g[37] | &p[54:37]&g[36] | &p[54:36]&g[35] | &p[54:35]&g[34] | &p[54:34]&g[33] | &p[54:33]&g[32] | &p[54:32]&g[31] | &p[54:31]&g[30] | &p[54:30]&g[29] | &p[54:29]&g[28] | &p[54:28]&g[27] | &p[54:27]&g[26] | &p[54:26]&g[25] | &p[54:25]&g[24] | &p[54:24]&g[23] | &p[54:23]&g[22] | &p[54:22]&g[21] | &p[54:21]&g[20] | &p[54:20]&g[19] | &p[54:19]&g[18] | &p[54:18]&g[17] | &p[54:17]&g[16] | &p[54:16]&g[15] | &p[54:15]&g[14] | &p[54:14]&g[13] | &p[54:13]&g[12] | &p[54:12]&g[11] | &p[54:11]&g[10] | &p[54:10]&g[9] | &p[54:9]&g[8] | &p[54:8]&g[7] | &p[54:7]&g[6] | &p[54:6]&g[5] | &p[54:5]&g[4] | &p[54:4]&g[3] | &p[54:3]&g[2] | &p[54:2]&g[1] | &p[54:1]&g[0] | &p[54:0]&c[0];
	assign c[56] = g[55] | &p[55:55]&g[54] | &p[55:54]&g[53] | &p[55:53]&g[52] | &p[55:52]&g[51] | &p[55:51]&g[50] | &p[55:50]&g[49] | &p[55:49]&g[48] | &p[55:48]&g[47] | &p[55:47]&g[46] | &p[55:46]&g[45] | &p[55:45]&g[44] | &p[55:44]&g[43] | &p[55:43]&g[42] | &p[55:42]&g[41] | &p[55:41]&g[40] | &p[55:40]&g[39] | &p[55:39]&g[38] | &p[55:38]&g[37] | &p[55:37]&g[36] | &p[55:36]&g[35] | &p[55:35]&g[34] | &p[55:34]&g[33] | &p[55:33]&g[32] | &p[55:32]&g[31] | &p[55:31]&g[30] | &p[55:30]&g[29] | &p[55:29]&g[28] | &p[55:28]&g[27] | &p[55:27]&g[26] | &p[55:26]&g[25] | &p[55:25]&g[24] | &p[55:24]&g[23] | &p[55:23]&g[22] | &p[55:22]&g[21] | &p[55:21]&g[20] | &p[55:20]&g[19] | &p[55:19]&g[18] | &p[55:18]&g[17] | &p[55:17]&g[16] | &p[55:16]&g[15] | &p[55:15]&g[14] | &p[55:14]&g[13] | &p[55:13]&g[12] | &p[55:12]&g[11] | &p[55:11]&g[10] | &p[55:10]&g[9] | &p[55:9]&g[8] | &p[55:8]&g[7] | &p[55:7]&g[6] | &p[55:6]&g[5] | &p[55:5]&g[4] | &p[55:4]&g[3] | &p[55:3]&g[2] | &p[55:2]&g[1] | &p[55:1]&g[0] | &p[55:0]&c[0];
	assign c[57] = g[56] | &p[56:56]&g[55] | &p[56:55]&g[54] | &p[56:54]&g[53] | &p[56:53]&g[52] | &p[56:52]&g[51] | &p[56:51]&g[50] | &p[56:50]&g[49] | &p[56:49]&g[48] | &p[56:48]&g[47] | &p[56:47]&g[46] | &p[56:46]&g[45] | &p[56:45]&g[44] | &p[56:44]&g[43] | &p[56:43]&g[42] | &p[56:42]&g[41] | &p[56:41]&g[40] | &p[56:40]&g[39] | &p[56:39]&g[38] | &p[56:38]&g[37] | &p[56:37]&g[36] | &p[56:36]&g[35] | &p[56:35]&g[34] | &p[56:34]&g[33] | &p[56:33]&g[32] | &p[56:32]&g[31] | &p[56:31]&g[30] | &p[56:30]&g[29] | &p[56:29]&g[28] | &p[56:28]&g[27] | &p[56:27]&g[26] | &p[56:26]&g[25] | &p[56:25]&g[24] | &p[56:24]&g[23] | &p[56:23]&g[22] | &p[56:22]&g[21] | &p[56:21]&g[20] | &p[56:20]&g[19] | &p[56:19]&g[18] | &p[56:18]&g[17] | &p[56:17]&g[16] | &p[56:16]&g[15] | &p[56:15]&g[14] | &p[56:14]&g[13] | &p[56:13]&g[12] | &p[56:12]&g[11] | &p[56:11]&g[10] | &p[56:10]&g[9] | &p[56:9]&g[8] | &p[56:8]&g[7] | &p[56:7]&g[6] | &p[56:6]&g[5] | &p[56:5]&g[4] | &p[56:4]&g[3] | &p[56:3]&g[2] | &p[56:2]&g[1] | &p[56:1]&g[0] | &p[56:0]&c[0];
	assign c[58] = g[57] | &p[57:57]&g[56] | &p[57:56]&g[55] | &p[57:55]&g[54] | &p[57:54]&g[53] | &p[57:53]&g[52] | &p[57:52]&g[51] | &p[57:51]&g[50] | &p[57:50]&g[49] | &p[57:49]&g[48] | &p[57:48]&g[47] | &p[57:47]&g[46] | &p[57:46]&g[45] | &p[57:45]&g[44] | &p[57:44]&g[43] | &p[57:43]&g[42] | &p[57:42]&g[41] | &p[57:41]&g[40] | &p[57:40]&g[39] | &p[57:39]&g[38] | &p[57:38]&g[37] | &p[57:37]&g[36] | &p[57:36]&g[35] | &p[57:35]&g[34] | &p[57:34]&g[33] | &p[57:33]&g[32] | &p[57:32]&g[31] | &p[57:31]&g[30] | &p[57:30]&g[29] | &p[57:29]&g[28] | &p[57:28]&g[27] | &p[57:27]&g[26] | &p[57:26]&g[25] | &p[57:25]&g[24] | &p[57:24]&g[23] | &p[57:23]&g[22] | &p[57:22]&g[21] | &p[57:21]&g[20] | &p[57:20]&g[19] | &p[57:19]&g[18] | &p[57:18]&g[17] | &p[57:17]&g[16] | &p[57:16]&g[15] | &p[57:15]&g[14] | &p[57:14]&g[13] | &p[57:13]&g[12] | &p[57:12]&g[11] | &p[57:11]&g[10] | &p[57:10]&g[9] | &p[57:9]&g[8] | &p[57:8]&g[7] | &p[57:7]&g[6] | &p[57:6]&g[5] | &p[57:5]&g[4] | &p[57:4]&g[3] | &p[57:3]&g[2] | &p[57:2]&g[1] | &p[57:1]&g[0] | &p[57:0]&c[0];
	assign c[59] = g[58] | &p[58:58]&g[57] | &p[58:57]&g[56] | &p[58:56]&g[55] | &p[58:55]&g[54] | &p[58:54]&g[53] | &p[58:53]&g[52] | &p[58:52]&g[51] | &p[58:51]&g[50] | &p[58:50]&g[49] | &p[58:49]&g[48] | &p[58:48]&g[47] | &p[58:47]&g[46] | &p[58:46]&g[45] | &p[58:45]&g[44] | &p[58:44]&g[43] | &p[58:43]&g[42] | &p[58:42]&g[41] | &p[58:41]&g[40] | &p[58:40]&g[39] | &p[58:39]&g[38] | &p[58:38]&g[37] | &p[58:37]&g[36] | &p[58:36]&g[35] | &p[58:35]&g[34] | &p[58:34]&g[33] | &p[58:33]&g[32] | &p[58:32]&g[31] | &p[58:31]&g[30] | &p[58:30]&g[29] | &p[58:29]&g[28] | &p[58:28]&g[27] | &p[58:27]&g[26] | &p[58:26]&g[25] | &p[58:25]&g[24] | &p[58:24]&g[23] | &p[58:23]&g[22] | &p[58:22]&g[21] | &p[58:21]&g[20] | &p[58:20]&g[19] | &p[58:19]&g[18] | &p[58:18]&g[17] | &p[58:17]&g[16] | &p[58:16]&g[15] | &p[58:15]&g[14] | &p[58:14]&g[13] | &p[58:13]&g[12] | &p[58:12]&g[11] | &p[58:11]&g[10] | &p[58:10]&g[9] | &p[58:9]&g[8] | &p[58:8]&g[7] | &p[58:7]&g[6] | &p[58:6]&g[5] | &p[58:5]&g[4] | &p[58:4]&g[3] | &p[58:3]&g[2] | &p[58:2]&g[1] | &p[58:1]&g[0] | &p[58:0]&c[0];
	assign c[60] = g[59] | &p[59:59]&g[58] | &p[59:58]&g[57] | &p[59:57]&g[56] | &p[59:56]&g[55] | &p[59:55]&g[54] | &p[59:54]&g[53] | &p[59:53]&g[52] | &p[59:52]&g[51] | &p[59:51]&g[50] | &p[59:50]&g[49] | &p[59:49]&g[48] | &p[59:48]&g[47] | &p[59:47]&g[46] | &p[59:46]&g[45] | &p[59:45]&g[44] | &p[59:44]&g[43] | &p[59:43]&g[42] | &p[59:42]&g[41] | &p[59:41]&g[40] | &p[59:40]&g[39] | &p[59:39]&g[38] | &p[59:38]&g[37] | &p[59:37]&g[36] | &p[59:36]&g[35] | &p[59:35]&g[34] | &p[59:34]&g[33] | &p[59:33]&g[32] | &p[59:32]&g[31] | &p[59:31]&g[30] | &p[59:30]&g[29] | &p[59:29]&g[28] | &p[59:28]&g[27] | &p[59:27]&g[26] | &p[59:26]&g[25] | &p[59:25]&g[24] | &p[59:24]&g[23] | &p[59:23]&g[22] | &p[59:22]&g[21] | &p[59:21]&g[20] | &p[59:20]&g[19] | &p[59:19]&g[18] | &p[59:18]&g[17] | &p[59:17]&g[16] | &p[59:16]&g[15] | &p[59:15]&g[14] | &p[59:14]&g[13] | &p[59:13]&g[12] | &p[59:12]&g[11] | &p[59:11]&g[10] | &p[59:10]&g[9] | &p[59:9]&g[8] | &p[59:8]&g[7] | &p[59:7]&g[6] | &p[59:6]&g[5] | &p[59:5]&g[4] | &p[59:4]&g[3] | &p[59:3]&g[2] | &p[59:2]&g[1] | &p[59:1]&g[0] | &p[59:0]&c[0];
	assign c[61] = g[60] | &p[60:60]&g[59] | &p[60:59]&g[58] | &p[60:58]&g[57] | &p[60:57]&g[56] | &p[60:56]&g[55] | &p[60:55]&g[54] | &p[60:54]&g[53] | &p[60:53]&g[52] | &p[60:52]&g[51] | &p[60:51]&g[50] | &p[60:50]&g[49] | &p[60:49]&g[48] | &p[60:48]&g[47] | &p[60:47]&g[46] | &p[60:46]&g[45] | &p[60:45]&g[44] | &p[60:44]&g[43] | &p[60:43]&g[42] | &p[60:42]&g[41] | &p[60:41]&g[40] | &p[60:40]&g[39] | &p[60:39]&g[38] | &p[60:38]&g[37] | &p[60:37]&g[36] | &p[60:36]&g[35] | &p[60:35]&g[34] | &p[60:34]&g[33] | &p[60:33]&g[32] | &p[60:32]&g[31] | &p[60:31]&g[30] | &p[60:30]&g[29] | &p[60:29]&g[28] | &p[60:28]&g[27] | &p[60:27]&g[26] | &p[60:26]&g[25] | &p[60:25]&g[24] | &p[60:24]&g[23] | &p[60:23]&g[22] | &p[60:22]&g[21] | &p[60:21]&g[20] | &p[60:20]&g[19] | &p[60:19]&g[18] | &p[60:18]&g[17] | &p[60:17]&g[16] | &p[60:16]&g[15] | &p[60:15]&g[14] | &p[60:14]&g[13] | &p[60:13]&g[12] | &p[60:12]&g[11] | &p[60:11]&g[10] | &p[60:10]&g[9] | &p[60:9]&g[8] | &p[60:8]&g[7] | &p[60:7]&g[6] | &p[60:6]&g[5] | &p[60:5]&g[4] | &p[60:4]&g[3] | &p[60:3]&g[2] | &p[60:2]&g[1] | &p[60:1]&g[0] | &p[60:0]&c[0];
	assign c[62] = g[61] | &p[61:61]&g[60] | &p[61:60]&g[59] | &p[61:59]&g[58] | &p[61:58]&g[57] | &p[61:57]&g[56] | &p[61:56]&g[55] | &p[61:55]&g[54] | &p[61:54]&g[53] | &p[61:53]&g[52] | &p[61:52]&g[51] | &p[61:51]&g[50] | &p[61:50]&g[49] | &p[61:49]&g[48] | &p[61:48]&g[47] | &p[61:47]&g[46] | &p[61:46]&g[45] | &p[61:45]&g[44] | &p[61:44]&g[43] | &p[61:43]&g[42] | &p[61:42]&g[41] | &p[61:41]&g[40] | &p[61:40]&g[39] | &p[61:39]&g[38] | &p[61:38]&g[37] | &p[61:37]&g[36] | &p[61:36]&g[35] | &p[61:35]&g[34] | &p[61:34]&g[33] | &p[61:33]&g[32] | &p[61:32]&g[31] | &p[61:31]&g[30] | &p[61:30]&g[29] | &p[61:29]&g[28] | &p[61:28]&g[27] | &p[61:27]&g[26] | &p[61:26]&g[25] | &p[61:25]&g[24] | &p[61:24]&g[23] | &p[61:23]&g[22] | &p[61:22]&g[21] | &p[61:21]&g[20] | &p[61:20]&g[19] | &p[61:19]&g[18] | &p[61:18]&g[17] | &p[61:17]&g[16] | &p[61:16]&g[15] | &p[61:15]&g[14] | &p[61:14]&g[13] | &p[61:13]&g[12] | &p[61:12]&g[11] | &p[61:11]&g[10] | &p[61:10]&g[9] | &p[61:9]&g[8] | &p[61:8]&g[7] | &p[61:7]&g[6] | &p[61:6]&g[5] | &p[61:5]&g[4] | &p[61:4]&g[3] | &p[61:3]&g[2] | &p[61:2]&g[1] | &p[61:1]&g[0] | &p[61:0]&c[0];
	assign c[63] = g[62] | &p[62:62]&g[61] | &p[62:61]&g[60] | &p[62:60]&g[59] | &p[62:59]&g[58] | &p[62:58]&g[57] | &p[62:57]&g[56] | &p[62:56]&g[55] | &p[62:55]&g[54] | &p[62:54]&g[53] | &p[62:53]&g[52] | &p[62:52]&g[51] | &p[62:51]&g[50] | &p[62:50]&g[49] | &p[62:49]&g[48] | &p[62:48]&g[47] | &p[62:47]&g[46] | &p[62:46]&g[45] | &p[62:45]&g[44] | &p[62:44]&g[43] | &p[62:43]&g[42] | &p[62:42]&g[41] | &p[62:41]&g[40] | &p[62:40]&g[39] | &p[62:39]&g[38] | &p[62:38]&g[37] | &p[62:37]&g[36] | &p[62:36]&g[35] | &p[62:35]&g[34] | &p[62:34]&g[33] | &p[62:33]&g[32] | &p[62:32]&g[31] | &p[62:31]&g[30] | &p[62:30]&g[29] | &p[62:29]&g[28] | &p[62:28]&g[27] | &p[62:27]&g[26] | &p[62:26]&g[25] | &p[62:25]&g[24] | &p[62:24]&g[23] | &p[62:23]&g[22] | &p[62:22]&g[21] | &p[62:21]&g[20] | &p[62:20]&g[19] | &p[62:19]&g[18] | &p[62:18]&g[17] | &p[62:17]&g[16] | &p[62:16]&g[15] | &p[62:15]&g[14] | &p[62:14]&g[13] | &p[62:13]&g[12] | &p[62:12]&g[11] | &p[62:11]&g[10] | &p[62:10]&g[9] | &p[62:9]&g[8] | &p[62:8]&g[7] | &p[62:7]&g[6] | &p[62:6]&g[5] | &p[62:5]&g[4] | &p[62:4]&g[3] | &p[62:3]&g[2] | &p[62:2]&g[1] | &p[62:1]&g[0] | &p[62:0]&c[0];
	assign c[64] = g[63] | &p[63:63]&g[62] | &p[63:62]&g[61] | &p[63:61]&g[60] | &p[63:60]&g[59] | &p[63:59]&g[58] | &p[63:58]&g[57] | &p[63:57]&g[56] | &p[63:56]&g[55] | &p[63:55]&g[54] | &p[63:54]&g[53] | &p[63:53]&g[52] | &p[63:52]&g[51] | &p[63:51]&g[50] | &p[63:50]&g[49] | &p[63:49]&g[48] | &p[63:48]&g[47] | &p[63:47]&g[46] | &p[63:46]&g[45] | &p[63:45]&g[44] | &p[63:44]&g[43] | &p[63:43]&g[42] | &p[63:42]&g[41] | &p[63:41]&g[40] | &p[63:40]&g[39] | &p[63:39]&g[38] | &p[63:38]&g[37] | &p[63:37]&g[36] | &p[63:36]&g[35] | &p[63:35]&g[34] | &p[63:34]&g[33] | &p[63:33]&g[32] | &p[63:32]&g[31] | &p[63:31]&g[30] | &p[63:30]&g[29] | &p[63:29]&g[28] | &p[63:28]&g[27] | &p[63:27]&g[26] | &p[63:26]&g[25] | &p[63:25]&g[24] | &p[63:24]&g[23] | &p[63:23]&g[22] | &p[63:22]&g[21] | &p[63:21]&g[20] | &p[63:20]&g[19] | &p[63:19]&g[18] | &p[63:18]&g[17] | &p[63:17]&g[16] | &p[63:16]&g[15] | &p[63:15]&g[14] | &p[63:14]&g[13] | &p[63:13]&g[12] | &p[63:12]&g[11] | &p[63:11]&g[10] | &p[63:10]&g[9] | &p[63:9]&g[8] | &p[63:8]&g[7] | &p[63:7]&g[6] | &p[63:6]&g[5] | &p[63:5]&g[4] | &p[63:4]&g[3] | &p[63:3]&g[2] | &p[63:2]&g[1] | &p[63:1]&g[0] | &p[63:0]&c[0];

	assign s = p^c[63:0];

	assign cOut = c[64];

endmodule
